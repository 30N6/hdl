library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library common_lib;
  use common_lib.common_pkg.all;

package eth_pkg is

end package eth_pkg;

package body eth_pkg is

end package body eth_pkg;
