library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library common_lib;
  use common_lib.common_pkg.all;
  use common_lib.math_pkg.all;

library dsp_lib;
  use dsp_lib.dsp_pkg.all;

entity channelized_dds_lut is
generic (
  DATA_WIDTH  : natural;
  LATENCY     : natural
);
port (
  Clk           : in  std_logic;

  Read_half     : in  std_logic;
  Read_index    : in  unsigned(DDS_SIN_LOOKUP_INDEX_WIDTH - 1 downto 0);

  Read_data     : out signed_array_t(1 downto 0)(DATA_WIDTH - 1 downto 0)
);
begin
  -- PSL default clock is rising_edge(Clk);
end entity channelized_dds_lut;

architecture rtl of channelized_dds_lut is

  constant LUT_WIDTH  : natural := 24;
  constant LUT_INIT   : std_logic_vector_array_t(2 ** DDS_SIN_LOOKUP_INDEX_WIDTH - 1 downto 0) :=
  (
       0 => "011111111111000000000000",    1 => "011111111111000000000110",    2 => "011111111111000000001101",    3 => "011111111111000000010011",    4 => "011111111111000000011001",    5 => "011111111111000000011111",    6 => "011111111111000000100110",    7 => "011111111111000000101100",
       8 => "011111111110000000110010",    9 => "011111111110000000111001",   10 => "011111111110000000111111",   11 => "011111111110000001000101",   12 => "011111111110000001001011",   13 => "011111111101000001010010",   14 => "011111111101000001011000",   15 => "011111111101000001011110",
      16 => "011111111101000001100100",   17 => "011111111100000001101011",   18 => "011111111100000001110001",   19 => "011111111100000001110111",   20 => "011111111011000001111110",   21 => "011111111011000010000100",   22 => "011111111010000010001010",   23 => "011111111010000010010000",
      24 => "011111111001000010010111",   25 => "011111111001000010011101",   26 => "011111111000000010100011",   27 => "011111111000000010101001",   28 => "011111110111000010110000",   29 => "011111110111000010110110",   30 => "011111110110000010111100",   31 => "011111110110000011000010",
      32 => "011111110101000011001001",   33 => "011111110101000011001111",   34 => "011111110100000011010101",   35 => "011111110011000011011011",   36 => "011111110011000011100010",   37 => "011111110010000011101000",   38 => "011111110001000011101110",   39 => "011111110000000011110100",
      40 => "011111110000000011111011",   41 => "011111101111000100000001",   42 => "011111101110000100000111",   43 => "011111101101000100001101",   44 => "011111101100000100010011",   45 => "011111101100000100011010",   46 => "011111101011000100100000",   47 => "011111101010000100100110",
      48 => "011111101001000100101100",   49 => "011111101000000100110011",   50 => "011111100111000100111001",   51 => "011111100110000100111111",   52 => "011111100101000101000101",   53 => "011111100100000101001011",   54 => "011111100011000101010010",   55 => "011111100010000101011000",
      56 => "011111100001000101011110",   57 => "011111100000000101100100",   58 => "011111011111000101101010",   59 => "011111011110000101110001",   60 => "011111011100000101110111",   61 => "011111011011000101111101",   62 => "011111011010000110000011",   63 => "011111011001000110001001",
      64 => "011111011000000110001111",   65 => "011111010110000110010110",   66 => "011111010101000110011100",   67 => "011111010100000110100010",   68 => "011111010011000110101000",   69 => "011111010001000110101110",   70 => "011111010000000110110100",   71 => "011111001111000110111010",
      72 => "011111001101000111000001",   73 => "011111001100000111000111",   74 => "011111001010000111001101",   75 => "011111001001000111010011",   76 => "011111001000000111011001",   77 => "011111000110000111011111",   78 => "011111000101000111100101",   79 => "011111000011000111101011",
      80 => "011111000010000111110001",   81 => "011111000000000111110111",   82 => "011110111111000111111110",   83 => "011110111101001000000100",   84 => "011110111011001000001010",   85 => "011110111010001000010000",   86 => "011110111000001000010110",   87 => "011110110111001000011100",
      88 => "011110110101001000100010",   89 => "011110110011001000101000",   90 => "011110110001001000101110",   91 => "011110110000001000110100",   92 => "011110101110001000111010",   93 => "011110101100001001000000",   94 => "011110101010001001000110",   95 => "011110101001001001001100",
      96 => "011110100111001001010010",   97 => "011110100101001001011000",   98 => "011110100011001001011110",   99 => "011110100001001001100100",  100 => "011110011111001001101010",  101 => "011110011110001001110000",  102 => "011110011100001001110110",  103 => "011110011010001001111100",
     104 => "011110011000001010000010",  105 => "011110010110001010001000",  106 => "011110010100001010001110",  107 => "011110010010001010010100",  108 => "011110010000001010011010",  109 => "011110001110001010100000",  110 => "011110001100001010100110",  111 => "011110001001001010101100",
     112 => "011110000111001010110010",  113 => "011110000101001010111000",  114 => "011110000011001010111101",  115 => "011110000001001011000011",  116 => "011101111111001011001001",  117 => "011101111101001011001111",  118 => "011101111010001011010101",  119 => "011101111000001011011011",
     120 => "011101110110001011100001",  121 => "011101110100001011100111",  122 => "011101110001001011101100",  123 => "011101101111001011110010",  124 => "011101101101001011111000",  125 => "011101101010001011111110",  126 => "011101101000001100000100",  127 => "011101100110001100001010",
     128 => "011101100011001100001111",  129 => "011101100001001100010101",  130 => "011101011110001100011011",  131 => "011101011100001100100001",  132 => "011101011001001100100111",  133 => "011101010111001100101100",  134 => "011101010100001100110010",  135 => "011101010010001100111000",
     136 => "011101001111001100111110",  137 => "011101001101001101000011",  138 => "011101001010001101001001",  139 => "011101001000001101001111",  140 => "011101000101001101010100",  141 => "011101000010001101011010",  142 => "011101000000001101100000",  143 => "011100111101001101100110",
     144 => "011100111010001101101011",  145 => "011100111000001101110001",  146 => "011100110101001101110111",  147 => "011100110010001101111100",  148 => "011100110000001110000010",  149 => "011100101101001110000111",  150 => "011100101010001110001101",  151 => "011100100111001110010011",
     152 => "011100100100001110011000",  153 => "011100100010001110011110",  154 => "011100011111001110100100",  155 => "011100011100001110101001",  156 => "011100011001001110101111",  157 => "011100010110001110110100",  158 => "011100010011001110111010",  159 => "011100010000001110111111",
     160 => "011100001101001111000101",  161 => "011100001010001111001010",  162 => "011100000111001111010000",  163 => "011100000100001111010110",  164 => "011100000001001111011011",  165 => "011011111110001111100001",  166 => "011011111011001111100110",  167 => "011011111000001111101011",
     168 => "011011110101001111110001",  169 => "011011110010001111110110",  170 => "011011101111001111111100",  171 => "011011101100010000000001",  172 => "011011101001010000000111",  173 => "011011100101010000001100",  174 => "011011100010010000010010",  175 => "011011011111010000010111",
     176 => "011011011100010000011100",  177 => "011011011001010000100010",  178 => "011011010101010000100111",  179 => "011011010010010000101100",  180 => "011011001111010000110010",  181 => "011011001011010000110111",  182 => "011011001000010000111101",  183 => "011011000101010001000010",
     184 => "011011000001010001000111",  185 => "011010111110010001001100",  186 => "011010111011010001010010",  187 => "011010110111010001010111",  188 => "011010110100010001011100",  189 => "011010110000010001100010",  190 => "011010101101010001100111",  191 => "011010101001010001101100",
     192 => "011010100110010001110001",  193 => "011010100011010001110110",  194 => "011010011111010001111100",  195 => "011010011011010010000001",  196 => "011010011000010010000110",  197 => "011010010100010010001011",  198 => "011010010001010010010000",  199 => "011010001101010010010110",
     200 => "011010001010010010011011",  201 => "011010000110010010100000",  202 => "011010000010010010100101",  203 => "011001111111010010101010",  204 => "011001111011010010101111",  205 => "011001110111010010110100",  206 => "011001110100010010111001",  207 => "011001110000010010111110",
     208 => "011001101100010011000011",  209 => "011001101000010011001000",  210 => "011001100101010011001101",  211 => "011001100001010011010010",  212 => "011001011101010011010111",  213 => "011001011001010011011100",  214 => "011001010101010011100001",  215 => "011001010010010011100110",
     216 => "011001001110010011101011",  217 => "011001001010010011110000",  218 => "011001000110010011110101",  219 => "011001000010010011111010",  220 => "011000111110010011111111",  221 => "011000111010010100000100",  222 => "011000110110010100001001",  223 => "011000110010010100001110",
     224 => "011000101110010100010011",  225 => "011000101010010100010111",  226 => "011000100110010100011100",  227 => "011000100010010100100001",  228 => "011000011110010100100110",  229 => "011000011010010100101011",  230 => "011000010110010100110000",  231 => "011000010010010100110100",
     232 => "011000001110010100111001",  233 => "011000001010010100111110",  234 => "011000000110010101000011",  235 => "011000000010010101000111",  236 => "010111111101010101001100",  237 => "010111111001010101010001",  238 => "010111110101010101010101",  239 => "010111110001010101011010",
     240 => "010111101101010101011111",  241 => "010111101001010101100011",  242 => "010111100100010101101000",  243 => "010111100000010101101101",  244 => "010111011100010101110001",  245 => "010111010111010101110110",  246 => "010111010011010101111010",  247 => "010111001111010101111111",
     248 => "010111001011010110000011",  249 => "010111000110010110001000",  250 => "010111000010010110001101",  251 => "010110111101010110010001",  252 => "010110111001010110010110",  253 => "010110110101010110011010",  254 => "010110110000010110011111",  255 => "010110101100010110100011",
     256 => "010110100111010110100111",  257 => "010110100011010110101100",  258 => "010110011111010110110000",  259 => "010110011010010110110101",  260 => "010110010110010110111001",  261 => "010110010001010110111101",  262 => "010110001101010111000010",  263 => "010110001000010111000110",
     264 => "010110000011010111001011",  265 => "010101111111010111001111",  266 => "010101111010010111010011",  267 => "010101110110010111010111",  268 => "010101110001010111011100",  269 => "010101101101010111100000",  270 => "010101101000010111100100",  271 => "010101100011010111101001",
     272 => "010101011111010111101101",  273 => "010101011010010111110001",  274 => "010101010101010111110101",  275 => "010101010001010111111001",  276 => "010101001100010111111101",  277 => "010101000111011000000010",  278 => "010101000011011000000110",  279 => "010100111110011000001010",
     280 => "010100111001011000001110",  281 => "010100110100011000010010",  282 => "010100110000011000010110",  283 => "010100101011011000011010",  284 => "010100100110011000011110",  285 => "010100100001011000100010",  286 => "010100011100011000100110",  287 => "010100010111011000101010",
     288 => "010100010011011000101110",  289 => "010100001110011000110010",  290 => "010100001001011000110110",  291 => "010100000100011000111010",  292 => "010011111111011000111110",  293 => "010011111010011001000010",  294 => "010011110101011001000110",  295 => "010011110000011001001010",
     296 => "010011101011011001001110",  297 => "010011100110011001010010",  298 => "010011100001011001010101",  299 => "010011011100011001011001",  300 => "010011010111011001011101",  301 => "010011010010011001100001",  302 => "010011001101011001100101",  303 => "010011001000011001101000",
     304 => "010011000011011001101100",  305 => "010010111110011001110000",  306 => "010010111001011001110100",  307 => "010010110100011001110111",  308 => "010010101111011001111011",  309 => "010010101010011001111111",  310 => "010010100101011010000010",  311 => "010010100000011010000110",
     312 => "010010011011011010001010",  313 => "010010010110011010001101",  314 => "010010010000011010010001",  315 => "010010001011011010010100",  316 => "010010000110011010011000",  317 => "010010000001011010011011",  318 => "010001111100011010011111",  319 => "010001110110011010100011",
     320 => "010001110001011010100110",  321 => "010001101100011010101001",  322 => "010001100111011010101101",  323 => "010001100010011010110000",  324 => "010001011100011010110100",  325 => "010001010111011010110111",  326 => "010001010010011010111011",  327 => "010001001100011010111110",
     328 => "010001000111011011000001",  329 => "010001000010011011000101",  330 => "010000111101011011001000",  331 => "010000110111011011001011",  332 => "010000110010011011001111",  333 => "010000101100011011010010",  334 => "010000100111011011010101",  335 => "010000100010011011011001",
     336 => "010000011100011011011100",  337 => "010000010111011011011111",  338 => "010000010010011011100010",  339 => "010000001100011011100101",  340 => "010000000111011011101001",  341 => "010000000001011011101100",  342 => "001111111100011011101111",  343 => "001111110110011011110010",
     344 => "001111110001011011110101",  345 => "001111101011011011111000",  346 => "001111100110011011111011",  347 => "001111100001011011111110",  348 => "001111011011011100000001",  349 => "001111010110011100000100",  350 => "001111010000011100000111",  351 => "001111001010011100001010",
     352 => "001111000101011100001101",  353 => "001110111111011100010000",  354 => "001110111010011100010011",  355 => "001110110100011100010110",  356 => "001110101111011100011001",  357 => "001110101001011100011100",  358 => "001110100100011100011111",  359 => "001110011110011100100010",
     360 => "001110011000011100100100",  361 => "001110010011011100100111",  362 => "001110001101011100101010",  363 => "001110000111011100101101",  364 => "001110000010011100110000",  365 => "001101111100011100110010",  366 => "001101110111011100110101",  367 => "001101110001011100111000",
     368 => "001101101011011100111010",  369 => "001101100110011100111101",  370 => "001101100000011101000000",  371 => "001101011010011101000010",  372 => "001101010100011101000101",  373 => "001101001111011101001000",  374 => "001101001001011101001010",  375 => "001101000011011101001101",
     376 => "001100111110011101001111",  377 => "001100111000011101010010",  378 => "001100110010011101010100",  379 => "001100101100011101010111",  380 => "001100100111011101011001",  381 => "001100100001011101011100",  382 => "001100011011011101011110",  383 => "001100010101011101100001",
     384 => "001100001111011101100011",  385 => "001100001010011101100110",  386 => "001100000100011101101000",  387 => "001011111110011101101010",  388 => "001011111000011101101101",  389 => "001011110010011101101111",  390 => "001011101100011101110001",  391 => "001011100111011101110100",
     392 => "001011100001011101110110",  393 => "001011011011011101111000",  394 => "001011010101011101111010",  395 => "001011001111011101111101",  396 => "001011001001011101111111",  397 => "001011000011011110000001",  398 => "001010111101011110000011",  399 => "001010111000011110000101",
     400 => "001010110010011110000111",  401 => "001010101100011110001001",  402 => "001010100110011110001100",  403 => "001010100000011110001110",  404 => "001010011010011110010000",  405 => "001010010100011110010010",  406 => "001010001110011110010100",  407 => "001010001000011110010110",
     408 => "001010000010011110011000",  409 => "001001111100011110011010",  410 => "001001110110011110011100",  411 => "001001110000011110011110",  412 => "001001101010011110011111",  413 => "001001100100011110100001",  414 => "001001011110011110100011",  415 => "001001011000011110100101",
     416 => "001001010010011110100111",  417 => "001001001100011110101001",  418 => "001001000110011110101010",  419 => "001001000000011110101100",  420 => "001000111010011110101110",  421 => "001000110100011110110000",  422 => "001000101110011110110001",  423 => "001000101000011110110011",
     424 => "001000100010011110110101",  425 => "001000011100011110110111",  426 => "001000010110011110111000",  427 => "001000010000011110111010",  428 => "001000001010011110111011",  429 => "001000000100011110111101",  430 => "000111111110011110111111",  431 => "000111110111011111000000",
     432 => "000111110001011111000010",  433 => "000111101011011111000011",  434 => "000111100101011111000101",  435 => "000111011111011111000110",  436 => "000111011001011111001000",  437 => "000111010011011111001001",  438 => "000111001101011111001010",  439 => "000111000111011111001100",
     440 => "000111000001011111001101",  441 => "000110111010011111001111",  442 => "000110110100011111010000",  443 => "000110101110011111010001",  444 => "000110101000011111010011",  445 => "000110100010011111010100",  446 => "000110011100011111010101",  447 => "000110010110011111010110",
     448 => "000110001111011111011000",  449 => "000110001001011111011001",  450 => "000110000011011111011010",  451 => "000101111101011111011011",  452 => "000101110111011111011100",  453 => "000101110001011111011110",  454 => "000101101010011111011111",  455 => "000101100100011111100000",
     456 => "000101011110011111100001",  457 => "000101011000011111100010",  458 => "000101010010011111100011",  459 => "000101001011011111100100",  460 => "000101000101011111100101",  461 => "000100111111011111100110",  462 => "000100111001011111100111",  463 => "000100110011011111101000",
     464 => "000100101100011111101001",  465 => "000100100110011111101010",  466 => "000100100000011111101011",  467 => "000100011010011111101100",  468 => "000100010011011111101100",  469 => "000100001101011111101101",  470 => "000100000111011111101110",  471 => "000100000001011111101111",
     472 => "000011111011011111110000",  473 => "000011110100011111110000",  474 => "000011101110011111110001",  475 => "000011101000011111110010",  476 => "000011100010011111110011",  477 => "000011011011011111110011",  478 => "000011010101011111110100",  479 => "000011001111011111110101",
     480 => "000011001001011111110101",  481 => "000011000010011111110110",  482 => "000010111100011111110110",  483 => "000010110110011111110111",  484 => "000010110000011111110111",  485 => "000010101001011111111000",  486 => "000010100011011111111000",  487 => "000010011101011111111001",
     488 => "000010010111011111111001",  489 => "000010010000011111111010",  490 => "000010001010011111111010",  491 => "000010000100011111111011",  492 => "000001111110011111111011",  493 => "000001110111011111111100",  494 => "000001110001011111111100",  495 => "000001101011011111111100",
     496 => "000001100100011111111101",  497 => "000001011110011111111101",  498 => "000001011000011111111101",  499 => "000001010010011111111101",  500 => "000001001011011111111110",  501 => "000001000101011111111110",  502 => "000000111111011111111110",  503 => "000000111001011111111110",
     504 => "000000110010011111111110",  505 => "000000101100011111111111",  506 => "000000100110011111111111",  507 => "000000011111011111111111",  508 => "000000011001011111111111",  509 => "000000010011011111111111",  510 => "000000001101011111111111",  511 => "000000000110011111111111",
     512 => "000000000000011111111111",  513 => "111111111010011111111111",  514 => "111111110011011111111111",  515 => "111111101101011111111111",  516 => "111111100111011111111111",  517 => "111111100001011111111111",  518 => "111111011010011111111111",  519 => "111111010100011111111111",
     520 => "111111001110011111111110",  521 => "111111000111011111111110",  522 => "111111000001011111111110",  523 => "111110111011011111111110",  524 => "111110110101011111111110",  525 => "111110101110011111111101",  526 => "111110101000011111111101",  527 => "111110100010011111111101",
     528 => "111110011100011111111101",  529 => "111110010101011111111100",  530 => "111110001111011111111100",  531 => "111110001001011111111100",  532 => "111110000010011111111011",  533 => "111101111100011111111011",  534 => "111101110110011111111010",  535 => "111101110000011111111010",
     536 => "111101101001011111111001",  537 => "111101100011011111111001",  538 => "111101011101011111111000",  539 => "111101010111011111111000",  540 => "111101010000011111110111",  541 => "111101001010011111110111",  542 => "111101000100011111110110",  543 => "111100111110011111110110",
     544 => "111100110111011111110101",  545 => "111100110001011111110101",  546 => "111100101011011111110100",  547 => "111100100101011111110011",  548 => "111100011110011111110011",  549 => "111100011000011111110010",  550 => "111100010010011111110001",  551 => "111100001100011111110000",
     552 => "111100000101011111110000",  553 => "111011111111011111101111",  554 => "111011111001011111101110",  555 => "111011110011011111101101",  556 => "111011101101011111101100",  557 => "111011100110011111101100",  558 => "111011100000011111101011",  559 => "111011011010011111101010",
     560 => "111011010100011111101001",  561 => "111011001101011111101000",  562 => "111011000111011111100111",  563 => "111011000001011111100110",  564 => "111010111011011111100101",  565 => "111010110101011111100100",  566 => "111010101110011111100011",  567 => "111010101000011111100010",
     568 => "111010100010011111100001",  569 => "111010011100011111100000",  570 => "111010010110011111011111",  571 => "111010001111011111011110",  572 => "111010001001011111011100",  573 => "111010000011011111011011",  574 => "111001111101011111011010",  575 => "111001110111011111011001",
     576 => "111001110001011111011000",  577 => "111001101010011111010110",  578 => "111001100100011111010101",  579 => "111001011110011111010100",  580 => "111001011000011111010011",  581 => "111001010010011111010001",  582 => "111001001100011111010000",  583 => "111001000110011111001111",
     584 => "111000111111011111001101",  585 => "111000111001011111001100",  586 => "111000110011011111001010",  587 => "111000101101011111001001",  588 => "111000100111011111001000",  589 => "111000100001011111000110",  590 => "111000011011011111000101",  591 => "111000010101011111000011",
     592 => "111000001111011111000010",  593 => "111000001001011111000000",  594 => "111000000010011110111111",  595 => "110111111100011110111101",  596 => "110111110110011110111011",  597 => "110111110000011110111010",  598 => "110111101010011110111000",  599 => "110111100100011110110111",
     600 => "110111011110011110110101",  601 => "110111011000011110110011",  602 => "110111010010011110110001",  603 => "110111001100011110110000",  604 => "110111000110011110101110",  605 => "110111000000011110101100",  606 => "110110111010011110101010",  607 => "110110110100011110101001",
     608 => "110110101110011110100111",  609 => "110110101000011110100101",  610 => "110110100010011110100011",  611 => "110110011100011110100001",  612 => "110110010110011110011111",  613 => "110110010000011110011110",  614 => "110110001010011110011100",  615 => "110110000100011110011010",
     616 => "110101111110011110011000",  617 => "110101111000011110010110",  618 => "110101110010011110010100",  619 => "110101101100011110010010",  620 => "110101100110011110010000",  621 => "110101100000011110001110",  622 => "110101011010011110001100",  623 => "110101010100011110001001",
     624 => "110101001110011110000111",  625 => "110101001000011110000101",  626 => "110101000011011110000011",  627 => "110100111101011110000001",  628 => "110100110111011101111111",  629 => "110100110001011101111101",  630 => "110100101011011101111010",  631 => "110100100101011101111000",
     632 => "110100011111011101110110",  633 => "110100011001011101110100",  634 => "110100010100011101110001",  635 => "110100001110011101101111",  636 => "110100001000011101101101",  637 => "110100000010011101101010",  638 => "110011111100011101101000",  639 => "110011110110011101100110",
     640 => "110011110001011101100011",  641 => "110011101011011101100001",  642 => "110011100101011101011110",  643 => "110011011111011101011100",  644 => "110011011001011101011001",  645 => "110011010100011101010111",  646 => "110011001110011101010100",  647 => "110011001000011101010010",
     648 => "110011000010011101001111",  649 => "110010111101011101001101",  650 => "110010110111011101001010",  651 => "110010110001011101001000",  652 => "110010101100011101000101",  653 => "110010100110011101000010",  654 => "110010100000011101000000",  655 => "110010011010011100111101",
     656 => "110010010101011100111010",  657 => "110010001111011100111000",  658 => "110010001001011100110101",  659 => "110010000100011100110010",  660 => "110001111110011100110000",  661 => "110001111001011100101101",  662 => "110001110011011100101010",  663 => "110001101101011100100111",
     664 => "110001101000011100100100",  665 => "110001100010011100100010",  666 => "110001011100011100011111",  667 => "110001010111011100011100",  668 => "110001010001011100011001",  669 => "110001001100011100010110",  670 => "110001000110011100010011",  671 => "110001000001011100010000",
     672 => "110000111011011100001101",  673 => "110000110110011100001010",  674 => "110000110000011100000111",  675 => "110000101010011100000100",  676 => "110000100101011100000001",  677 => "110000011111011011111110",  678 => "110000011010011011111011",  679 => "110000010101011011111000",
     680 => "110000001111011011110101",  681 => "110000001010011011110010",  682 => "110000000100011011101111",  683 => "101111111111011011101100",  684 => "101111111001011011101001",  685 => "101111110100011011100101",  686 => "101111101110011011100010",  687 => "101111101001011011011111",
     688 => "101111100100011011011100",  689 => "101111011110011011011001",  690 => "101111011001011011010101",  691 => "101111010100011011010010",  692 => "101111001110011011001111",  693 => "101111001001011011001011",  694 => "101111000011011011001000",  695 => "101110111110011011000101",
     696 => "101110111001011011000001",  697 => "101110110100011010111110",  698 => "101110101110011010111011",  699 => "101110101001011010110111",  700 => "101110100100011010110100",  701 => "101110011110011010110000",  702 => "101110011001011010101101",  703 => "101110010100011010101001",
     704 => "101110001111011010100110",  705 => "101110001010011010100011",  706 => "101110000100011010011111",  707 => "101101111111011010011011",  708 => "101101111010011010011000",  709 => "101101110101011010010100",  710 => "101101110000011010010001",  711 => "101101101010011010001101",
     712 => "101101100101011010001010",  713 => "101101100000011010000110",  714 => "101101011011011010000010",  715 => "101101010110011001111111",  716 => "101101010001011001111011",  717 => "101101001100011001110111",  718 => "101101000111011001110100",  719 => "101101000010011001110000",
     720 => "101100111101011001101100",  721 => "101100111000011001101000",  722 => "101100110011011001100101",  723 => "101100101110011001100001",  724 => "101100101001011001011101",  725 => "101100100100011001011001",  726 => "101100011111011001010101",  727 => "101100011010011001010010",
     728 => "101100010101011001001110",  729 => "101100010000011001001010",  730 => "101100001011011001000110",  731 => "101100000110011001000010",  732 => "101100000001011000111110",  733 => "101011111100011000111010",  734 => "101011110111011000110110",  735 => "101011110010011000110010",
     736 => "101011101101011000101110",  737 => "101011101001011000101010",  738 => "101011100100011000100110",  739 => "101011011111011000100010",  740 => "101011011010011000011110",  741 => "101011010101011000011010",  742 => "101011010000011000010110",  743 => "101011001100011000010010",
     744 => "101011000111011000001110",  745 => "101011000010011000001010",  746 => "101010111101011000000110",  747 => "101010111001011000000010",  748 => "101010110100010111111101",  749 => "101010101111010111111001",  750 => "101010101011010111110101",  751 => "101010100110010111110001",
     752 => "101010100001010111101101",  753 => "101010011101010111101001",  754 => "101010011000010111100100",  755 => "101010010011010111100000",  756 => "101010001111010111011100",  757 => "101010001010010111010111",  758 => "101010000110010111010011",  759 => "101010000001010111001111",
     760 => "101001111101010111001011",  761 => "101001111000010111000110",  762 => "101001110011010111000010",  763 => "101001101111010110111101",  764 => "101001101010010110111001",  765 => "101001100110010110110101",  766 => "101001100001010110110000",  767 => "101001011101010110101100",
     768 => "101001011001010110100111",  769 => "101001010100010110100011",  770 => "101001010000010110011111",  771 => "101001001011010110011010",  772 => "101001000111010110010110",  773 => "101001000011010110010001",  774 => "101000111110010110001101",  775 => "101000111010010110001000",
     776 => "101000110101010110000011",  777 => "101000110001010101111111",  778 => "101000101101010101111010",  779 => "101000101001010101110110",  780 => "101000100100010101110001",  781 => "101000100000010101101101",  782 => "101000011100010101101000",  783 => "101000010111010101100011",
     784 => "101000010011010101011111",  785 => "101000001111010101011010",  786 => "101000001011010101010101",  787 => "101000000111010101010001",  788 => "101000000011010101001100",  789 => "100111111110010101000111",  790 => "100111111010010101000011",  791 => "100111110110010100111110",
     792 => "100111110010010100111001",  793 => "100111101110010100110100",  794 => "100111101010010100110000",  795 => "100111100110010100101011",  796 => "100111100010010100100110",  797 => "100111011110010100100001",  798 => "100111011010010100011100",  799 => "100111010110010100010111",
     800 => "100111010010010100010011",  801 => "100111001110010100001110",  802 => "100111001010010100001001",  803 => "100111000110010100000100",  804 => "100111000010010011111111",  805 => "100110111110010011111010",  806 => "100110111010010011110101",  807 => "100110110110010011110000",
     808 => "100110110010010011101011",  809 => "100110101110010011100110",  810 => "100110101011010011100001",  811 => "100110100111010011011100",  812 => "100110100011010011010111",  813 => "100110011111010011010010",  814 => "100110011011010011001101",  815 => "100110011000010011001000",
     816 => "100110010100010011000011",  817 => "100110010000010010111110",  818 => "100110001100010010111001",  819 => "100110001001010010110100",  820 => "100110000101010010101111",  821 => "100110000001010010101010",  822 => "100101111110010010100101",  823 => "100101111010010010100000",
     824 => "100101110110010010011011",  825 => "100101110011010010010110",  826 => "100101101111010010010000",  827 => "100101101100010010001011",  828 => "100101101000010010000110",  829 => "100101100101010010000001",  830 => "100101100001010001111100",  831 => "100101011101010001110110",
     832 => "100101011010010001110001",  833 => "100101010111010001101100",  834 => "100101010011010001100111",  835 => "100101010000010001100010",  836 => "100101001100010001011100",  837 => "100101001001010001010111",  838 => "100101000101010001010010",  839 => "100101000010010001001100",
     840 => "100100111111010001000111",  841 => "100100111011010001000010",  842 => "100100111000010000111101",  843 => "100100110101010000110111",  844 => "100100110001010000110010",  845 => "100100101110010000101100",  846 => "100100101011010000100111",  847 => "100100100111010000100010",
     848 => "100100100100010000011100",  849 => "100100100001010000010111",  850 => "100100011110010000010010",  851 => "100100011011010000001100",  852 => "100100010111010000000111",  853 => "100100010100010000000001",  854 => "100100010001001111111100",  855 => "100100001110001111110110",
     856 => "100100001011001111110001",  857 => "100100001000001111101011",  858 => "100100000101001111100110",  859 => "100100000010001111100001",  860 => "100011111111001111011011",  861 => "100011111100001111010110",  862 => "100011111001001111010000",  863 => "100011110110001111001010",
     864 => "100011110011001111000101",  865 => "100011110000001110111111",  866 => "100011101101001110111010",  867 => "100011101010001110110100",  868 => "100011100111001110101111",  869 => "100011100100001110101001",  870 => "100011100001001110100100",  871 => "100011011110001110011110",
     872 => "100011011100001110011000",  873 => "100011011001001110010011",  874 => "100011010110001110001101",  875 => "100011010011001110000111",  876 => "100011010000001110000010",  877 => "100011001110001101111100",  878 => "100011001011001101110111",  879 => "100011001000001101110001",
     880 => "100011000110001101101011",  881 => "100011000011001101100110",  882 => "100011000000001101100000",  883 => "100010111110001101011010",  884 => "100010111011001101010100",  885 => "100010111000001101001111",  886 => "100010110110001101001001",  887 => "100010110011001101000011",
     888 => "100010110001001100111110",  889 => "100010101110001100111000",  890 => "100010101100001100110010",  891 => "100010101001001100101100",  892 => "100010100111001100100111",  893 => "100010100100001100100001",  894 => "100010100010001100011011",  895 => "100010011111001100010101",
     896 => "100010011101001100001111",  897 => "100010011010001100001010",  898 => "100010011000001100000100",  899 => "100010010110001011111110",  900 => "100010010011001011111000",  901 => "100010010001001011110010",  902 => "100010001111001011101100",  903 => "100010001100001011100111",
     904 => "100010001010001011100001",  905 => "100010001000001011011011",  906 => "100010000110001011010101",  907 => "100010000011001011001111",  908 => "100010000001001011001001",  909 => "100001111111001011000011",  910 => "100001111101001010111101",  911 => "100001111011001010111000",
     912 => "100001111001001010110010",  913 => "100001110111001010101100",  914 => "100001110100001010100110",  915 => "100001110010001010100000",  916 => "100001110000001010011010",  917 => "100001101110001010010100",  918 => "100001101100001010001110",  919 => "100001101010001010001000",
     920 => "100001101000001010000010",  921 => "100001100110001001111100",  922 => "100001100100001001110110",  923 => "100001100010001001110000",  924 => "100001100001001001101010",  925 => "100001011111001001100100",  926 => "100001011101001001011110",  927 => "100001011011001001011000",
     928 => "100001011001001001010010",  929 => "100001010111001001001100",  930 => "100001010110001001000110",  931 => "100001010100001001000000",  932 => "100001010010001000111010",  933 => "100001010000001000110100",  934 => "100001001111001000101110",  935 => "100001001101001000101000",
     936 => "100001001011001000100010",  937 => "100001001001001000011100",  938 => "100001001000001000010110",  939 => "100001000110001000010000",  940 => "100001000101001000001010",  941 => "100001000011001000000100",  942 => "100001000001000111111110",  943 => "100001000000000111110111",
     944 => "100000111110000111110001",  945 => "100000111101000111101011",  946 => "100000111011000111100101",  947 => "100000111010000111011111",  948 => "100000111000000111011001",  949 => "100000110111000111010011",  950 => "100000110110000111001101",  951 => "100000110100000111000111",
     952 => "100000110011000111000001",  953 => "100000110001000110111010",  954 => "100000110000000110110100",  955 => "100000101111000110101110",  956 => "100000101101000110101000",  957 => "100000101100000110100010",  958 => "100000101011000110011100",  959 => "100000101010000110010110",
     960 => "100000101000000110001111",  961 => "100000100111000110001001",  962 => "100000100110000110000011",  963 => "100000100101000101111101",  964 => "100000100100000101110111",  965 => "100000100010000101110001",  966 => "100000100001000101101010",  967 => "100000100000000101100100",
     968 => "100000011111000101011110",  969 => "100000011110000101011000",  970 => "100000011101000101010010",  971 => "100000011100000101001011",  972 => "100000011011000101000101",  973 => "100000011010000100111111",  974 => "100000011001000100111001",  975 => "100000011000000100110011",
     976 => "100000010111000100101100",  977 => "100000010110000100100110",  978 => "100000010101000100100000",  979 => "100000010100000100011010",  980 => "100000010100000100010011",  981 => "100000010011000100001101",  982 => "100000010010000100000111",  983 => "100000010001000100000001",
     984 => "100000010000000011111011",  985 => "100000010000000011110100",  986 => "100000001111000011101110",  987 => "100000001110000011101000",  988 => "100000001101000011100010",  989 => "100000001101000011011011",  990 => "100000001100000011010101",  991 => "100000001011000011001111",
     992 => "100000001011000011001001",  993 => "100000001010000011000010",  994 => "100000001010000010111100",  995 => "100000001001000010110110",  996 => "100000001001000010110000",  997 => "100000001000000010101001",  998 => "100000001000000010100011",  999 => "100000000111000010011101",
    1000 => "100000000111000010010111", 1001 => "100000000110000010010000", 1002 => "100000000110000010001010", 1003 => "100000000101000010000100", 1004 => "100000000101000001111110", 1005 => "100000000100000001110111", 1006 => "100000000100000001110001", 1007 => "100000000100000001101011",
    1008 => "100000000011000001100100", 1009 => "100000000011000001011110", 1010 => "100000000011000001011000", 1011 => "100000000011000001010010", 1012 => "100000000010000001001011", 1013 => "100000000010000001000101", 1014 => "100000000010000000111111", 1015 => "100000000010000000111001",
    1016 => "100000000010000000110010", 1017 => "100000000001000000101100", 1018 => "100000000001000000100110", 1019 => "100000000001000000011111", 1020 => "100000000001000000011001", 1021 => "100000000001000000010011", 1022 => "100000000001000000001101", 1023 => "100000000001000000000110"
  );

  signal m_lut          : std_logic_vector_array_t(2 ** DDS_SIN_LOOKUP_INDEX_WIDTH - 1 downto 0)(LUT_WIDTH - 1 downto 0) := LUT_INIT;

  signal r0_read_half   : std_logic;
  signal r0_read_data   : std_logic_vector(LUT_WIDTH - 1 downto 0);

  signal r1_read_half   : std_logic;
  signal r1_read_data   : std_logic_vector(LUT_WIDTH - 1 downto 0);
  signal w1_data_i      : signed(LUT_WIDTH/2 - 1 downto 0);
  signal w1_data_q      : signed(LUT_WIDTH/2 - 1 downto 0);
  signal w1_data_i_inv  : signed(LUT_WIDTH/2 - 1 downto 0);
  signal w1_data_q_inv  : signed(LUT_WIDTH/2 - 1 downto 0);

begin

  assert (LATENCY = 3)
    report "LATENCY expected to be 3"
    severity failure;

  assert (DATA_WIDTH = LUT_WIDTH/2)
    report "DATA_WIDTH must be = LUT_WIDTH/2, otherwise max negative->invert behavior is not guaranteed"
    severity failure;

  process(Clk)
  begin
    if rising_edge(Clk) then
      r0_read_half <= Read_half;
      r0_read_data <= m_lut(to_integer(Read_index));
    end if;
  end process;

  process(Clk)
  begin
    if rising_edge(Clk) then
      r1_read_half <= r0_read_half;
      r1_read_data <= r0_read_data;
    end if;
  end process;

  (w1_data_q, w1_data_i) <= signed(r1_read_data);
  w1_data_i_inv <= -w1_data_i;
  w1_data_q_inv <= -w1_data_q;

  -- PSL underflow_i : assert always (w1_data_i(LUT_WIDTH/2 - 1) = '1') -> (or_reduce(w1_data_i(LUT_WIDTH/2 - 2 downto 0)) = '1');
  -- PSL underflow_q : assert always (w1_data_q(LUT_WIDTH/2 - 1) = '1') -> (or_reduce(w1_data_q(LUT_WIDTH/2 - 2 downto 0)) = '1');

  process(Clk)
  begin
    if rising_edge(Clk) then
      if (r1_read_half = '0') then
        Read_data(0) <= w1_data_i(LUT_WIDTH/2 - 1 downto (LUT_WIDTH/2 - DATA_WIDTH));
        Read_data(1) <= w1_data_q(LUT_WIDTH/2 - 1 downto (LUT_WIDTH/2 - DATA_WIDTH));
      else
        Read_data(0) <= w1_data_i_inv(LUT_WIDTH/2 - 1 downto (LUT_WIDTH/2 - DATA_WIDTH));
        Read_data(1) <= w1_data_q_inv(LUT_WIDTH/2 - 1 downto (LUT_WIDTH/2 - DATA_WIDTH));
      end if;
    end if;
  end process;

end architecture rtl;
