library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library common_lib;
  use common_lib.common_pkg.all;

package esm_pkg is

  constant ESM_CONTROL_MAGIC_NUM                        : std_logic_vector(31 downto 0) := "45534D43";
  constant ESM_REPORT_MAGIC_NUM                         : std_logic_vector(31 downto 0) := "45534D52";

  constant ESM_MODULE_ID_WIDTH                          : natural := 2;
  constant ESM_MESSAGE_TYPE_WIDTH                       : natural := 8;

  constant ESM_MODULE_ID_CONTROL                        : unsigned(ESM_MODULE_ID_WIDTH - 1 downto 0) := "00";
  constant ESM_MODULE_ID_DWELL                          : unsigned(ESM_MODULE_ID_WIDTH - 1 downto 0) := "01";
  constant ESM_MODULE_ID_PDW                            : unsigned(ESM_MODULE_ID_WIDTH - 1 downto 0) := "10";

  constant ESM_CONTROL_MESSAGE_TYPE_ENABLE              : unsigned(ESM_MESSAGE_TYPE_WIDTH - 1 downto 0) := x"00";
  constant ESM_CONTROL_MESSAGE_TYPE_DWELL_ENTRY         : unsigned(ESM_MESSAGE_TYPE_WIDTH - 1 downto 0) := x"01";
  constant ESM_CONTROL_MESSAGE_TYPE_DWELL_PROGRAM       : unsigned(ESM_MESSAGE_TYPE_WIDTH - 1 downto 0) := x"02";
  constant ESM_CONTROL_MESSAGE_TYPE_PDW_SETUP           : unsigned(ESM_MESSAGE_TYPE_WIDTH - 1 downto 0) := x"03";  --TODO: unused?

  constant ESM_REPORT_MESSAGE_TYPE_DWELL_COMPLETE_INFO  : unsigned(ESM_MESSAGE_TYPE_WIDTH - 1 downto 0) := x"10";
  constant ESM_REPORT_MESSAGE_TYPE_DWELL_COMPLETE_STATS : unsigned(ESM_MESSAGE_TYPE_WIDTH - 1 downto 0) := x"10";
  constant ESM_REPORT_MESSAGE_TYPE_PDW                  : unsigned(ESM_MESSAGE_TYPE_WIDTH - 1 downto 0) := x"20";

  constant ESM_NUM_CHANNELS_NARROW                      : natural := 64;
  constant ESM_NUM_CHANNELS_WIDE                        : natural := 8;
  constant ESM_CHANNEL_INDEX_WIDTH                      : natural := clog2(ESM_NUM_CHANNELS_WIDE);

  constant ESM_NUM_FAST_LOCK_PROFILES                   : natural := 8;
  constant ESM_FAST_LOCK_PROFILE_INDEX_WIDTH            : natural := clog2(ESM_NUM_FAST_LOCK_PROFILES);
  constant ESM_NUM_DWELL_ENTRIES                        : natural := 32;
  constant ESM_DWELL_ENTRY_INDEX_WIDTH                  : natural := clog2(ESM_NUM_DWELL_ENTRIES);
  constant ESM_NUM_DWELL_INSTRUCTIONS                   : natural := 32;
  constant ESM_DWELL_INSTRUCTION_INDEX_WIDTH            : natural := clog2(ESM_NUM_DWELL_INSTRUCTIONS);

  --type esm_common_header_t is record
  --  magic_num                 : std_logic_vector(31 downto 0);
  --  sequence_num              : unsigned(31 downto 0);
  --  module_id                 : unsigned(ESM_MODULE_ID_WIDTH - 1 downto 0);
  --  message_type              : unsigned(ESM_MESSAGE_TYPE_WIDTH - 1 downto 0);
  --end record;

  --type esm_message_enable_t is record
  --  header                    : esm_common_header_t;
  --  reset                     : std_logic;
  --  enable_channelizer        : std_logic_vector(1 downto 0);
  --  enable_pdw                : std_logic_vector(1 downto 0);
  --end record;

  type esm_dwell_metadata_t is record
    tag                       : unsigned(15 downto 0);
    frequency                 : unsigned(15 downto 0);
    duration                  : unsigned(31 downto 0);
    gain                      : unsigned(6 downto 0);
    fast_lock_profile         : unsigned(ESM_FAST_LOCK_PROFILE_INDEX_WIDTH - 1 downto 0);
    threshold_narrow          : unsigned(15 downto 0);
    threshold_wide            : unsigned(15 downto 0);
    channel_mask_narrow       : std_logic_vector(ESM_NUM_CHANNELS_NARROW - 1 downto 0);
    channel_mask_wide         : std_logic_vector(ESM_NUM_CHANNELS_WIDE - 1 downto 0);
  end record;

  type esm_dwell_metadata_array_t is array (natural range <>) of esm_dwell_metadata_t;

  constant ESM_DWELL_METADATA_PACKED_WIDTH : natural := 184;
  --type esm_dwell_metadata_packed_t is record
  --  tag                       : unsigned(15 downto 0);
  --  frequency                 : unsigned(15 downto 0);
  --  duration                  : unsigned(31 downto 0);
  --  gain                      : unsigned(7 downto 0);
  --  fast_lock_profile         : unsigned(7 downto 0);
  --  threshold_narrow          : unsigned(15 downto 0);
  --  threshold_wide            : unsigned(15 downto 0);
  --  channel_mask_narrow       : std_logic_vector(63 downto 0);
  --  channel_mask_wide         : std_logic_vector(7 downto 0);
  --end record;

  type esm_message_dwell_entry_t is record
    entry_index               : unsigned(ESM_DWELL_ENTRY_INDEX_WIDTH - 1 downto 0);
    entry_data                : esm_dwell_metadata_t;
  end record;

  constant ESM_MESSAGE_DWELL_ENTRY_PACKED_WIDTH : natural := 8 + ESM_DWELL_METADATA_PACKED_WIDTH;
  --type esm_message_dwell_entry_packed_t is record
  --  entry_index               : unsigned(7 downto 0);
  --  entry_data                : esm_dwell_metadata_packed_t;
  --end record;

  type esm_dwell_instruction_t is record
    valid                     : std_logic;
    global_counter_check      : std_logic;
    global_counter_dec        : std_logic;
    repeat_count              : unsigned(3 downto 0);
    entry_index               : unsigned(ESM_DWELL_ENTRY_INDEX_WIDTH - 1 downto 0);
    next_instruction_index    : unsigned(ESM_DWELL_INSTRUCTION_INDEX_WIDTH - 1 downto 0);
  end record;

  constant ESM_DWELL_INSTRUCTION_PACKED_WIDTH : natural := 32;
  --type esm_message_dwell_instruction_packed_t is record
  --  flags                     : std_logic_vector(7 downto 0);
  --  repeat_count              : unsigned(7 downto 0);
  --  entry_index               : unsigned(7 downto 0);
  --  next_instruction_index    : unsigned(7 downto 0);
  --end record;

  type esm_dwell_instruction_array_t is array (natural range <>) of esm_dwell_instruction_t;

  --type esm_message_dwell_program_t is record
  --  --header                    : esm_common_header_t;
  --  enable_program            : std_logic;
  --  enable_delayed_start      : std_logic;
  --  global_counter_init       : unsigned(31 downto 0);
  --  delayed_start_time        : unsigned(63 downto 0);
  --  instructions              : esm_dwell_instruction_array_t(ESM_NUM_DWELL_INSTRUCTIONS - 1 downto 0);
  --end record;

  type esm_message_dwell_program_header_t is record
    enable_program            : std_logic;
    enable_delayed_start      : std_logic;
    global_counter_init       : unsigned(31 downto 0);
    delayed_start_time        : unsigned(63 downto 0);
  end record;

  constant ESM_MESSAGE_DWELL_PROGRAM_HEADER_PACKED_WIDTH : natural := 128;
  --type esm_message_dwell_program_header_packed_t is record
  --  --header                    : esm_common_header_t;
  --  enable_program            : std_logic_vector(7 downto 0);
  --  enable_delayed_start      : std_logic_vector(7 downto 0);
  --  padding                   : std_logic_vector(15 downto 0);
  --  global_counter_init       : unsigned(31 downto 0);
  --  delayed_start_time        : unsigned(63 downto 0);
  --  --instructions              : esm_dwell_instruction_array_packed_t(ESM_NUM_DWELL_INSTRUCTIONS - 1 downto 0);
  --end record;

  type esm_message_dwell_complete_info_t is record
    header                    : esm_common_header_t;
    dwell_sequence_num        : unsigned(31 downto 0);
    metadata                  : esm_dwell_metadata_t;

    num_samples               : unsigned(31 downto 0);
    ts_dwell_start            : unsigned(63 downto 0);
    ts_pll_locked             : unsigned(63 downto 0);
    ts_dwell_end              : unsigned(63 downto 0);
  end record;

  type esm_message_dwell_complete_stats_t is record
    header                    : esm_common_header_t;
    dwell_sequence_num        : unsigned(31 downto 0);
    metadata                  : esm_dwell_metadata_t;

    channel_start_index       : unsigned(ESM_CHANNEL_INDEX_WIDTH - 1 downto 0);
    channel_amplitude         : unsigned_array_t(ESM_NUM_CHANNELS_WIDE/2 - 1 downto 0)(31 downto 0);
  end record;

  type esm_message_pdw_t is record
    header                    : esm_common_header_t;
    pdw_sequence_num          : unsigned(31 downto 0);
    dwell_sequence_num        : unsigned(31 downto 0);
    dwell_metadata            : esm_dwell_metadata_t;
    pulse_channel             : unsigned(ESM_CHANNEL_INDEX_WIDTH - 1 downto 0);
    pulse_threshold           : unsigned(31 downto 0);
    pulse_amplitude           : unsigned(31 downto 0);
    pulse_duration            : unsigned(31 downto 0);  --TODO: early termination flag?
    pulse_frequency           : unsigned(31 downto 0);  --TODO: IFM module
    pulse_start_time          : unsigned(63 downto 0);
    raw_samples               : std_logic_vector_array_t(40 downto 0)(31 downto 0); --TODO: increase to max
  end record;

  type esm_config_data_t is record
    valid                     : std_logic;
    first                     : std_logic;
    last                      : std_logic;
    data                      : std_logic_vector(31 downto 0);
    module_id                 : unsigned(ESM_MODULE_ID_WIDTH - 1 downto 0);
    message_type              : unsigned(ESM_MESSAGE_TYPE_WIDTH - 1 downto 0);
  end record;

  function unpack(v : std_logic_vector) return esm_dwell_metadata_t;
  function unpack(v : std_logic_vector) return esm_message_dwell_entry_t;
  function unpack(v : std_logic_vector) return esm_message_dwell_program_header_t;
  function unpack(v : std_logic_vector) return esm_dwell_instruction_t;

end package esm_pkg;

package body esm_pkg is

  function unpack(v : std_logic_vector) return esm_dwell_metadata_t is
    variable r : esm_dwell_metadata_t;
  begin
    assert (v'length = ESM_DWELL_METADATA_PACKED_WIDTH)
      report "Unexpected length"
      severity failure;

    r.tag                 := v(15 downto 0);
    r.frequency           := v(31 downto 16);
    r.duration            := v(63 downto 32);
    r.gain                := v(70 downto 64);
    r.fast_lock_profile   := v(74 downto 72);
    r.threshold_narrow    := v(95 downto 80);
    r.threshold_wide      := v(111 downto 96);
    r.channel_mask_narrow := v(175 downto 112);
    r.channel_mask_wide   := v(183 downto 176);
    return r;
  end function;

  function unpack(v : std_logic_vector) return esm_message_dwell_entry_t is
    variable r : esm_message_dwell_entry_t;
  begin
    assert (v'length = ESM_MESSAGE_DWELL_ENTRY_PACKED_WIDTH)
      report "Unexpected length"
      severity failure;

    r.entry_index   := v(ESM_DWELL_ENTRY_INDEX_WIDTH - 1 downto 0);
    r.entry_data    := unpack(v(8 + ESM_DWELL_METADATA_PACKED_WIDTH - 1 downto 8));
    return r;
  end function;

  function unpack(v : std_logic_vector) return esm_message_dwell_program_header_t is
    variable r : esm_message_dwell_program_header_t;
  begin
    assert (v'length = ESM_MESSAGE_DWELL_PROGRAM_HEADER_PACKED_WIDTH)
      report "Unexpected length"
      severity failure;

    r.enable_program        := v(0);
    r.enable_delayed_start  := v(8);
    r.global_counter_init   := v(63 downto 32);
    r.delayed_start_time    := v(127 downto 64);
    return r;
  end function;

  function unpack(v : std_logic_vector) return esm_dwell_instruction_t is
    variable r : esm_dwell_instruction_t;
  begin
    assert (v'length = ESM_DWELL_INSTRUCTION_PACKED_WIDTH)
      report "Unexpected length"
      severity failure;

    r.valid                   := v(0);
    r.global_counter_check    := v(1);
    r.global_counter_dec      := v(2);
    r.repeat_count            := v(11 downto 8);
    r.entry_index             := v(20 downto 16);
    r.next_instruction_index  := v(28 downto 24);
    return r;
  end function;

end package body esm_pkg;
