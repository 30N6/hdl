library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library common_lib;
  use common_lib.common_pkg.all;
  use common_lib.math_pkg.all;

library dsp_lib;
  use dsp_lib.dsp_pkg.all;

entity synthesizer_16 is
generic (
  INPUT_DATA_WIDTH  : natural;
  OUTPUT_DATA_WIDTH : natural
);
port (
  Clk                       : in  std_logic;
  Rst                       : in  std_logic;

  Input_ctrl                : in  channelizer_control_t;
  Input_data                : in  signed_array_t(1 downto 0)(INPUT_DATA_WIDTH - 1 downto 0);

  Output_valid              : out std_logic;
  Output_data               : out signed_array_t(1 downto 0)(OUTPUT_DATA_WIDTH - 1 downto 0);

  Error_stretcher_overflow  : out std_logic;
  Error_stretcher_underflow : out std_logic;
  Error_filter_overflow     : out std_logic;
  Error_mux_input_overflow  : out std_logic;
  Error_mux_fifo_overflow   : out std_logic;
  Error_mux_fifo_underflow  : out std_logic
);
end entity synthesizer_16;

architecture rtl of synthesizer_16 is

  constant NUM_CHANNELS : natural := 16;
  constant NUM_COEFS    : natural := 192;
  constant COEF_WIDTH   : natural := 20;
  constant COEF_DATA    : signed_array_t(NUM_COEFS - 1 downto 0)(COEF_WIDTH - 1 downto 0) := (
      0 => "00000000000000000011",   1 => "00000000000000000000",   2 => "11111111111111111001",   3 => "11111111111111101110",   4 => "11111111111111011110",   5 => "11111111111111001000",   6 => "11111111111110101101",   7 => "11111111111110001100",
      8 => "11111111111101101000",   9 => "11111111111101000011",  10 => "11111111111100100000",  11 => "11111111111100000101",  12 => "11111111111011110101",  13 => "11111111111011110110",  14 => "11111111111100001111",  15 => "11111111111101000101",
     16 => "11111111111110011110",  17 => "00000000000000011101",  18 => "00000000000011000011",  19 => "00000000000110010010",  20 => "00000000001010000100",  21 => "00000000001110010011",  22 => "00000000010010110011",  23 => "00000000010111010110",
     24 => "00000000011011101001",  25 => "00000000011111010101",  26 => "00000000100010000010",  27 => "00000000100011010110",  28 => "00000000100010110111",  29 => "00000000100000001100",  30 => "00000000011011000001",  31 => "00000000010011001000",
     32 => "00000000001000011000",  33 => "11111111111010110011",  34 => "11111111101010101000",  35 => "11111111011000010000",  36 => "11111111000100010011",  37 => "11111110101111100100",  38 => "11111110011011000011",  39 => "11111110000111111100",
     40 => "11111101110111100010",  41 => "11111101101011001101",  42 => "11111101100100010100",  43 => "11111101100100001101",  44 => "11111101101100000000",  45 => "11111101111100101000",  46 => "11111110010110101100",  47 => "11111110111010010110",
     48 => "11111111100111010101",  49 => "00000000011100110011",  50 => "00000001011001010111",  51 => "00000010011011000011",  52 => "00000011011111011000",  53 => "00000100100011010100",  54 => "00000101100011011100",  55 => "00000110011100000100",
     56 => "00000111001001010101",  57 => "00000111100111011010",  58 => "00000111110010101100",  59 => "00000111101000000001",  60 => "00000111000100110110",  61 => "00000110000111011110",  62 => "00000100101111001101",  63 => "00000010111100100010",
     64 => "00000000110001010010",  65 => "11111110010000100110",  66 => "11111011011111000011",  67 => "11111000100010100011",  68 => "11110101100010010010",  69 => "11110010100110011110",  70 => "11101111111000010001",  71 => "11101101100001010101",
     72 => "11101011101011100110",  73 => "11101010100000111001",  74 => "11101010001010100010",  75 => "11101010110000111000",  76 => "11101100011011000011",  77 => "11101111001110011111",  78 => "11110011001110100111",  79 => "11111000011100101010",
     80 => "11111110110111011001",  81 => "00000110011011000000",  82 => "00001111000001001001",  83 => "00011000100000111110",  84 => "00100010101111010110",  85 => "00101101011111000011",  86 => "00111000100001001110",  87 => "01000011100101101100",
     88 => "01001110011011100011",  89 => "01011000110001101100",  90 => "01100010010111010010",  91 => "01101010111100011010",  92 => "01110010010010100011",  93 => "01111000001101001001",  94 => "01111100100001111011",  95 => "01111111001001011001",
     96 => "01111111111110111111",  97 => "01111111000001010010",  98 => "01111100010010000011",  99 => "01110111110110001011", 100 => "01110001110101011100", 101 => "01101010011010010111", 102 => "01100001110001101101", 103 => "01011000001010000111",
    104 => "01001101110011100101", 105 => "01000010111110111010", 106 => "00110111111101001011", 107 => "00101100111111001000", 108 => "00100010010100101111", 109 => "00011000001100100111", 110 => "00001110110011101100", 111 => "00000110010100110101",
    112 => "11111110111000100011", 113 => "11111000100100111010", 114 => "11110011011101011001", 115 => "11101111100010111111", 116 => "11101100110100010010", 117 => "11101011001101101011", 118 => "11101010101001100110", 119 => "11101011000000111011",
    120 => "11101100001011010001", 121 => "11101101111111011001", 122 => "11110000010011100110", 123 => "11110010111110001000", 124 => "11110101110101011111", 125 => "11111000110000110001", 126 => "11111011100111111110", 127 => "11111110010100001010",
    128 => "00000000101111101001", 129 => "00000010110110000100", 130 => "00000100100100011101", 131 => "00000101111001001000", 132 => "00000110110011101111", 133 => "00000111010100111111", 134 => "00000111011110101001", 135 => "00000111010011001101",
    136 => "00000110110101110100", 137 => "00000110001001111101", 138 => "00000101010011010111", 139 => "00000100010101110000", 140 => "00000011010100101100", 141 => "00000010010011011011", 142 => "00000001010100110110", 143 => "00000000011011010011",
    144 => "11111111101000101001", 145 => "11111110111110001010", 146 => "11111110011100100111", 147 => "11111110000100001101", 148 => "11111101110100110001", 149 => "11111101101101101011", 150 => "11111101101110000010", 151 => "11111101110100101110",
    152 => "11111110000000100000", 153 => "11111110010000000010", 154 => "11111110100010000010", 155 => "11111110110101010001", 156 => "11111111001000101001", 157 => "11111111011011001110", 158 => "11111111101100010001", 159 => "11111111111011001101",
    160 => "00000000000111101100", 161 => "00000000010001100010", 162 => "00000000011000101110", 163 => "00000000011101011000", 164 => "00000000011111101110", 165 => "00000000100000000101", 166 => "00000000011110110011", 167 => "00000000011100010001",
    168 => "00000000011000110111", 169 => "00000000010100111100", 170 => "00000000010000110011", 171 => "00000000001100101111", 172 => "00000000001000111011", 173 => "00000000000101100011", 174 => "00000000000010101100", 175 => "00000000000000011001",
    176 => "11111111111110101010", 177 => "11111111111101011110", 178 => "11111111111100110001", 179 => "11111111111100011101", 180 => "11111111111100011101", 181 => "11111111111100101100", 182 => "11111111111101000101", 183 => "11111111111101100100",
    184 => "11111111111110000100", 185 => "11111111111110100011", 186 => "11111111111110111110", 187 => "11111111111111010101", 188 => "11111111111111100110", 189 => "11111111111111110011", 190 => "11111111111111111011", 191 => "00000000000000000000"
  );

begin

  i_synthesizer : entity dsp_lib.synthesizer_common
  generic map (
    INPUT_DATA_WIDTH  => INPUT_DATA_WIDTH,
    OUTPUT_DATA_WIDTH => OUTPUT_DATA_WIDTH,
    NUM_CHANNELS      => NUM_CHANNELS,
    NUM_COEFS         => NUM_COEFS,
    COEF_WIDTH        => COEF_WIDTH,
    COEF_DATA         => COEF_DATA
  )
  port map (
    Clk                       => Clk,
    Rst                       => Rst,


    Input_ctrl                => Input_ctrl,
    Input_data                => Input_data,

    Output_valid              => Output_valid,
    Output_data               => Output_data,

    Error_stretcher_overflow  => Error_stretcher_overflow,
    Error_stretcher_underflow => Error_stretcher_underflow,
    Error_filter_overflow     => Error_filter_overflow,
    Error_mux_input_overflow  => Error_mux_input_overflow,
    Error_mux_fifo_overflow   => Error_mux_fifo_overflow,
    Error_mux_fifo_underflow  => Error_mux_fifo_underflow
  );

end architecture rtl;
