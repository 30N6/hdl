library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library common_lib;
  use common_lib.common_pkg.all;
  use common_lib.math_pkg.all;

library dsp_lib;
  use dsp_lib.dsp_pkg.all;

entity channelized_dds_lut is
generic (
  DATA_WIDTH  : natural;
  LATENCY     : natural
);
port (
  Clk           : in  std_logic;

  Read_half     : in  std_logic;
  Read_index    : in  unsigned(DDS_SIN_LOOKUP_INDEX_WIDTH - 1 downto 0);

  Read_data     : out signed_array_t(1 downto 0)(DATA_WIDTH - 1 downto 0)
);
begin
  -- PSL default clock is rising_edge(Clk);
end entity channelized_dds_lut;

architecture rtl of channelized_dds_lut is

  constant LUT_WIDTH  : natural := 32;
  constant LUT_INIT   : std_logic_vector_array_t(2 ** DDS_SIN_LOOKUP_INDEX_WIDTH - 1 downto 0) :=
  (
       0 => "01111111111111110000000000000000",    1 => "01111111111111110000000001100101",    2 => "01111111111111100000000011001001",    3 => "01111111111111100000000100101110",    4 => "01111111111111010000000110010010",    5 => "01111111111110110000000111110111",    6 => "01111111111110010000001001011011",    7 => "01111111111101110000001011000000",
       8 => "01111111111101010000001100100100",    9 => "01111111111100110000001110001001",   10 => "01111111111100000000001111101101",   11 => "01111111111011000000010001010010",   12 => "01111111111010010000010010110110",   13 => "01111111111001010000010100011011",   14 => "01111111111000010000010101111111",   15 => "01111111110111000000010111100011",
      16 => "01111111110110000000011001001000",   17 => "01111111110100100000011010101100",   18 => "01111111110011010000011100010001",   19 => "01111111110001110000011101110101",   20 => "01111111110000010000011111011001",   21 => "01111111101110110000100000111110",   22 => "01111111101101000000100010100010",   23 => "01111111101011010000100100000110",
      24 => "01111111101001100000100101101010",   25 => "01111111100111110000100111001111",   26 => "01111111100101110000101000110011",   27 => "01111111100011110000101010010111",   28 => "01111111100001100000101011111011",   29 => "01111111011111010000101101011111",   30 => "01111111011101000000101111000100",   31 => "01111111011010110000110000101000",
      32 => "01111111011000010000110010001100",   33 => "01111111010101110000110011110000",   34 => "01111111010011010000110101010100",   35 => "01111111010000100000110110111000",   36 => "01111111001101110000111000011100",   37 => "01111111001011000000111010000000",   38 => "01111111001000010000111011100011",   39 => "01111111000101010000111101000111",
      40 => "01111111000010010000111110101011",   41 => "01111110111111000001000000001111",   42 => "01111110111011110001000001110010",   43 => "01111110111000100001000011010110",   44 => "01111110110101010001000100111010",   45 => "01111110110001110001000110011101",   46 => "01111110101110010001001000000001",   47 => "01111110101010110001001001100100",
      48 => "01111110100111000001001011001000",   49 => "01111110100011010001001100101011",   50 => "01111110011111100001001110001111",   51 => "01111110011011110001001111110010",   52 => "01111110010111110001010001010101",   53 => "01111110010011110001010010111001",   54 => "01111110001111100001010100011100",   55 => "01111110001011100001010101111111",
      56 => "01111110000111010001010111100010",   57 => "01111110000010110001011001000101",   58 => "01111101111110100001011010101000",   59 => "01111101111010000001011100001011",   60 => "01111101110101010001011101101110",   61 => "01111101110000110001011111010000",   62 => "01111101101100000001100000110011",   63 => "01111101100111010001100010010110",
      64 => "01111101100010010001100011111001",   65 => "01111101011101100001100101011011",   66 => "01111101011000100001100110111110",   67 => "01111101010011010001101000100000",   68 => "01111101001110010001101010000010",   69 => "01111101001001000001101011100101",   70 => "01111101000011100001101101000111",   71 => "01111100111110010001101110101001",
      72 => "01111100111000110001110000001011",   73 => "01111100110011010001110001101101",   74 => "01111100101101100001110011001111",   75 => "01111100100111110001110100110001",   76 => "01111100100010000001110110010011",   77 => "01111100011100010001110111110101",   78 => "01111100010110010001111001010111",   79 => "01111100010000010001111010111000",
      80 => "01111100001010010001111100011010",   81 => "01111100000100000001111101111011",   82 => "01111011111110000001111111011101",   83 => "01111011110111100010000000111110",   84 => "01111011110001010010000010011111",   85 => "01111011101010110010000100000000",   86 => "01111011100100010010000101100001",   87 => "01111011011101110010000111000010",
      88 => "01111011010111000010001000100011",   89 => "01111011010000010010001010000100",   90 => "01111011001001100010001011100101",   91 => "01111011000010100010001101000110",   92 => "01111010111011100010001110100110",   93 => "01111010110100100010010000000111",   94 => "01111010101101100010010001100111",   95 => "01111010100110010010010011001000",
      96 => "01111010011111000010010100101000",   97 => "01111010010111110010010110001000",   98 => "01111010010000010010010111101000",   99 => "01111010001000110010011001001000",  100 => "01111010000001010010011010101000",  101 => "01111001111001100010011100001000",  102 => "01111001110010000010011101100111",  103 => "01111001101010010010011111000111",
     104 => "01111001100010010010100000100110",  105 => "01111001011010100010100010000110",  106 => "01111001010010100010100011100101",  107 => "01111001001010010010100101000100",  108 => "01111001000010010010100110100011",  109 => "01111000111010000010101000000010",  110 => "01111000110001110010101001100001",  111 => "01111000101001010010101011000000",
     112 => "01111000100001000010101100011111",  113 => "01111000011000100010101101111101",  114 => "01111000001111110010101111011100",  115 => "01111000000111010010110000111010",  116 => "01110111111110100010110010011001",  117 => "01110111110101110010110011110111",  118 => "01110111101100110010110101010101",  119 => "01110111100011110010110110110011",
     120 => "01110111011010110010111000010001",  121 => "01110111010001110010111001101110",  122 => "01110111001000100010111011001100",  123 => "01110110111111100010111100101010",  124 => "01110110110110000010111110000111",  125 => "01110110101100110010111111100100",  126 => "01110110100011010011000001000001",  127 => "01110110011001110011000010011110",
     128 => "01110110010000010011000011111011",  129 => "01110110000110100011000101011000",  130 => "01110101111100110011000110110101",  131 => "01110101110011000011001000010001",  132 => "01110101101001010011001001101110",  133 => "01110101011111010011001011001010",  134 => "01110101010101010011001100100110",  135 => "01110101001011010011001110000011",
     136 => "01110101000001000011001111011111",  137 => "01110100110110110011010000111010",  138 => "01110100101100100011010010010110",  139 => "01110100100010000011010011110010",  140 => "01110100010111110011010101001101",  141 => "01110100001101010011010110101000",  142 => "01110100000010100011011000000100",  143 => "01110011111000000011011001011111",
     144 => "01110011101101010011011010111010",  145 => "01110011100010100011011100010101",  146 => "01110011010111100011011101101111",  147 => "01110011001100110011011111001010",  148 => "01110011000001110011100000100100",  149 => "01110010110110110011100001111110",  150 => "01110010101011100011100011011001",  151 => "01110010100000010011100100110011",
     152 => "01110010010101000011100110001100",  153 => "01110010001001110011100111100110",  154 => "01110001111110010011101001000000",  155 => "01110001110010110011101010011001",  156 => "01110001100111010011101011110010",  157 => "01110001011011110011101101001100",  158 => "01110001010000000011101110100101",  159 => "01110001000100010011101111111110",
     160 => "01110000111000100011110001010110",  161 => "01110000101100100011110010101111",  162 => "01110000100000110011110100000111",  163 => "01110000010100110011110101100000",  164 => "01110000001000100011110110111000",  165 => "01101111111100100011111000010000",  166 => "01101111110000010011111001101000",  167 => "01101111100100000011111010111111",
     168 => "01101111010111100011111100010111",  169 => "01101111001011000011111101101110",  170 => "01101110111110110011111111000101",  171 => "01101110110010000100000000011101",  172 => "01101110100101100100000001110011",  173 => "01101110011000110100000011001010",  174 => "01101110001100000100000100100001",  175 => "01101101111111010100000101110111",
     176 => "01101101110010010100000111001110",  177 => "01101101100101010100001000100100",  178 => "01101101011000010100001001111010",  179 => "01101101001011010100001011010000",  180 => "01101100111110000100001100100101",  181 => "01101100110000110100001101111011",  182 => "01101100100011100100001111010000",  183 => "01101100010110010100010000100101",
     184 => "01101100001000110100010001111010",  185 => "01101011111011010100010011001111",  186 => "01101011101101110100010100100100",  187 => "01101011100000010100010101111000",  188 => "01101011010010100100010111001101",  189 => "01101011000100110100011000100001",  190 => "01101010110111000100011001110101",  191 => "01101010101001000100011011001001",
     192 => "01101010011011010100011100011100",  193 => "01101010001101010100011101110000",  194 => "01101001111111010100011111000011",  195 => "01101001110001000100100000010110",  196 => "01101001100010110100100001101001",  197 => "01101001010100100100100010111100",  198 => "01101001000110010100100100001111",  199 => "01101000111000000100100101100001",
     200 => "01101000101001100100100110110100",  201 => "01101000011011000100101000000110",  202 => "01101000001100100100101001011000",  203 => "01100111111101110100101010101001",  204 => "01100111101111000100101011111011",  205 => "01100111100000010100101101001100",  206 => "01100111010001100100101110011101",  207 => "01100111000010100100101111101110",
     208 => "01100110110011110100110000111111",  209 => "01100110100100110100110010010000",  210 => "01100110010101100100110011100000",  211 => "01100110000110100100110100110001",  212 => "01100101110111010100110110000001",  213 => "01100101101000000100110111010001",  214 => "01100101011000110100111000100000",  215 => "01100101001001010100111001110000",
     216 => "01100100111010000100111010111111",  217 => "01100100101010100100111100001110",  218 => "01100100011011000100111101011101",  219 => "01100100001011010100111110101100",  220 => "01100011111011100100111111111011",  221 => "01100011101011110101000001001001",  222 => "01100011011100000101000010010111",  223 => "01100011001100010101000011100101",
     224 => "01100010111100010101000100110011",  225 => "01100010101100010101000110000001",  226 => "01100010011100010101000111001110",  227 => "01100010001100010101001000011011",  228 => "01100001111100000101001001101000",  229 => "01100001101011110101001010110101",  230 => "01100001011011100101001100000010",  231 => "01100001001011010101001101001110",
     232 => "01100000111010110101001110011011",  233 => "01100000101010100101001111100111",  234 => "01100000011010000101010000110010",  235 => "01100000001001010101010001111110",  236 => "01011111111000110101010011001001",  237 => "01011111101000000101010100010101",  238 => "01011111010111010101010101100000",  239 => "01011111000110100101010110101010",
     240 => "01011110110101110101010111110101",  241 => "01011110100100110101011000111111",  242 => "01011110010011110101011010001010",  243 => "01011110000010110101011011010011",  244 => "01011101110001110101011100011101",  245 => "01011101100000100101011101100111",  246 => "01011101001111100101011110110000",  247 => "01011100111110010101011111111001",
     248 => "01011100101100110101100001000010",  249 => "01011100011011100101100010001011",  250 => "01011100001010000101100011010011",  251 => "01011011111000100101100100011100",  252 => "01011011100111000101100101100100",  253 => "01011011010101100101100110101100",  254 => "01011011000011110101100111110011",  255 => "01011010110010010101101000111011",
     256 => "01011010100000100101101010000010",  257 => "01011010001110110101101011001001",  258 => "01011001111100110101101100001111",  259 => "01011001101011000101101101010110",  260 => "01011001011001000101101110011100",  261 => "01011001000111000101101111100010",  262 => "01011000110100110101110000101000",  263 => "01011000100010110101110001101110",
     264 => "01011000010000100101110010110011",  265 => "01010111111110010101110011111001",  266 => "01010111101100000101110100111110",  267 => "01010111011001110101110110000010",  268 => "01010111000111010101110111000111",  269 => "01010110110100110101111000001011",  270 => "01010110100010100101111001001111",  271 => "01010110001111110101111010010011",
     272 => "01010101111101010101111011010111",  273 => "01010101101010100101111100011010",  274 => "01010101011000000101111101011101",  275 => "01010101000101010101111110100000",  276 => "01010100110010010101111111100011",  277 => "01010100011111100110000000100101",  278 => "01010100001100100110000001101000",  279 => "01010011111001110110000010101010",
     280 => "01010011100110110110000011101011",  281 => "01010011010011100110000100101101",  282 => "01010011000000100110000101101110",  283 => "01010010101101010110000110101111",  284 => "01010010011010000110000111110000",  285 => "01010010000110110110001000110001",  286 => "01010001110011100110001001110001",  287 => "01010001100000010110001010110001",
     288 => "01010001001100110110001011110001",  289 => "01010000111001010110001100110001",  290 => "01010000100101110110001101110000",  291 => "01010000010010010110001110101111",  292 => "01001111111110110110001111101110",  293 => "01001111101011000110010000101101",  294 => "01001111010111010110010001101100",  295 => "01001111000011100110010010101010",
     296 => "01001110101111110110010011101000",  297 => "01001110011100000110010100100101",  298 => "01001110001000000110010101100011",  299 => "01001101110100010110010110100000",  300 => "01001101100000010110010111011101",  301 => "01001101001100010110011000011010",  302 => "01001100111000000110011001010110",  303 => "01001100100100000110011010010011",
     304 => "01001100001111110110011011001111",  305 => "01001011111011100110011100001010",  306 => "01001011100111010110011101000110",  307 => "01001011010011000110011110000001",  308 => "01001010111110110110011110111100",  309 => "01001010101010010110011111110111",  310 => "01001010010110000110100000110010",  311 => "01001010000001100110100001101100",
     312 => "01001001101101000110100010100110",  313 => "01001001011000010110100011100000",  314 => "01001001000011110110100100011001",  315 => "01001000101111000110100101010010",  316 => "01001000011010010110100110001011",  317 => "01001000000101100110100111000100",  318 => "01000111110000110110100111111101",  319 => "01000111011100000110101000110101",
     320 => "01000111000111000110101001101101",  321 => "01000110110010010110101010100100",  322 => "01000110011101010110101011011100",  323 => "01000110001000010110101100010011",  324 => "01000101110011010110101101001010",  325 => "01000101011110000110101110000001",  326 => "01000101001001000110101110110111",  327 => "01000100110011110110101111101101",
     328 => "01000100011110100110110000100011",  329 => "01000100001001010110110001011001",  330 => "01000011110100000110110010001110",  331 => "01000011011110110110110011000011",  332 => "01000011001001010110110011111000",  333 => "01000010110100000110110100101101",  334 => "01000010011110100110110101100001",  335 => "01000010001001000110110110010101",
     336 => "01000001110011100110110111001001",  337 => "01000001011101110110110111111101",  338 => "01000001001000010110111000110000",  339 => "01000000110010100110111001100011",  340 => "01000000011100110110111010010110",  341 => "01000000000111010110111011001000",  342 => "00111111110001010110111011111011",  343 => "00111111011011100110111100101100",
     344 => "00111111000101110110111101011110",  345 => "00111110101111110110111110010000",  346 => "00111110011010000110111111000001",  347 => "00111110000100000110111111110010",  348 => "00111101101110000111000000100010",  349 => "00111101011000000111000001010011",  350 => "00111101000001110111000010000011",  351 => "00111100101011110111000010110010",
     352 => "00111100010101100111000011100010",  353 => "00111011111111100111000100010001",  354 => "00111011101001010111000101000000",  355 => "00111011010011000111000101101111",  356 => "00111010111100100111000110011101",  357 => "00111010100110010111000111001011",  358 => "00111010010000000111000111111001",  359 => "00111001111001100111001000100111",
     360 => "00111001100011000111001001010100",  361 => "00111001001100110111001010000001",  362 => "00111000110110010111001010101110",  363 => "00111000011111100111001011011011",  364 => "00111000001001000111001100000111",  365 => "00110111110010100111001100110011",  366 => "00110111011011110111001101011110",  367 => "00110111000101010111001110001010",
     368 => "00110110101110100111001110110101",  369 => "00110110010111110111001111100000",  370 => "00110110000001000111010000001010",  371 => "00110101101010000111010000110101",  372 => "00110101010011010111010001011111",  373 => "00110100111100100111010010001000",  374 => "00110100100101100111010010110010",  375 => "00110100001110100111010011011011",
     376 => "00110011110111110111010100000100",  377 => "00110011100000110111010100101101",  378 => "00110011001001100111010101010101",  379 => "00110010110010100111010101111101",  380 => "00110010011011100111010110100101",  381 => "00110010000100010111010111001100",  382 => "00110001101101010111010111110011",  383 => "00110001010110000111011000011010",
     384 => "00110000111110110111011001000001",  385 => "00110000100111100111011001100111",  386 => "00110000010000010111011010001101",  387 => "00101111111001000111011010110011",  388 => "00101111100001110111011011011000",  389 => "00101111001010100111011011111110",  390 => "00101110110011000111011100100010",  391 => "00101110011011100111011101000111",
     392 => "00101110000100010111011101101011",  393 => "00101101101100110111011110001111",  394 => "00101101010101010111011110110011",  395 => "00101100111101110111011111010111",  396 => "00101100100110010111011111111010",  397 => "00101100001110100111100000011101",  398 => "00101011110111000111100000111111",  399 => "00101011011111010111100001100010",
     400 => "00101011000111110111100010000100",  401 => "00101010110000000111100010100101",  402 => "00101010011000010111100011000111",  403 => "00101010000000100111100011101000",  404 => "00101001101000110111100100001001",  405 => "00101001010001000111100100101001",  406 => "00101000111001010111100101001010",  407 => "00101000100001100111100101101010",
     408 => "00101000001001100111100110001001",  409 => "00100111110001110111100110101001",  410 => "00100111011001110111100111001000",  411 => "00100111000010000111100111100110",  412 => "00100110101010000111101000000101",  413 => "00100110010010000111101000100011",  414 => "00100101111010000111101001000001",  415 => "00100101100010000111101001011111",
     416 => "00100101001010000111101001111100",  417 => "00100100110010000111101010011001",  418 => "00100100011001110111101010110110",  419 => "00100100000001110111101011010010",  420 => "00100011101001100111101011101110",  421 => "00100011010001100111101100001010",  422 => "00100010111001010111101100100110",  423 => "00100010100001000111101101000001",
     424 => "00100010001000110111101101011100",  425 => "00100001110000100111101101110111",  426 => "00100001011000010111101110010001",  427 => "00100001000000000111101110101011",  428 => "00100000100111110111101111000101",  429 => "00100000001111100111101111011110",  430 => "00011111110111010111101111111000",  431 => "00011111011110110111110000010000",
     432 => "00011111000110100111110000101001",  433 => "00011110101110000111110001000001",  434 => "00011110010101110111110001011001",  435 => "00011101111101010111110001110001",  436 => "00011101100100110111110010001000",  437 => "00011101001100010111110010011111",  438 => "00011100110011110111110010110110",  439 => "00011100011011010111110011001101",
     440 => "00011100000010110111110011100011",  441 => "00011011101010010111110011111001",  442 => "00011011010001110111110100001110",  443 => "00011010111001010111110100100100",  444 => "00011010100000100111110100111001",  445 => "00011010001000000111110101001101",  446 => "00011001101111100111110101100010",  447 => "00011001010110110111110101110110",
     448 => "00011000111110010111110110001001",  449 => "00011000100101100111110110011101",  450 => "00011000001100110111110110110000",  451 => "00010111110100000111110111000011",  452 => "00010111011011100111110111010101",  453 => "00010111000010110111110111101000",  454 => "00010110101010000111110111111010",  455 => "00010110010001010111111000001011",
     456 => "00010101111000100111111000011101",  457 => "00010101011111110111111000101110",  458 => "00010101000111000111111000111110",  459 => "00010100101110010111111001001111",  460 => "00010100010101010111111001011111",  461 => "00010011111100100111111001101111",  462 => "00010011100011110111111001111110",  463 => "00010011001010110111111010001101",
     464 => "00010010110010000111111010011100",  465 => "00010010011001000111111010101011",  466 => "00010010000000010111111010111001",  467 => "00010001100111010111111011000111",  468 => "00010001001110100111111011010101",  469 => "00010000110101100111111011100010",  470 => "00010000011100100111111011101111",  471 => "00010000000011110111111011111100",
     472 => "00001111101010110111111100001001",  473 => "00001111010001110111111100010101",  474 => "00001110111000110111111100100001",  475 => "00001110100000000111111100101100",  476 => "00001110000111000111111100110111",  477 => "00001101101110000111111101000010",  478 => "00001101010101000111111101001101",  479 => "00001100111100000111111101010111",
     480 => "00001100100011000111111101100001",  481 => "00001100001010000111111101101011",  482 => "00001011110001000111111101110100",  483 => "00001011010111110111111101111101",  484 => "00001010111110110111111110000110",  485 => "00001010100101110111111110001111",  486 => "00001010001100110111111110010111",  487 => "00001001110011110111111110011111",
     488 => "00001001011010100111111110100110",  489 => "00001001000001100111111110101101",  490 => "00001000101000100111111110110100",  491 => "00001000001111100111111110111011",  492 => "00000111110110010111111111000001",  493 => "00000111011101010111111111000111",  494 => "00000111000100010111111111001101",  495 => "00000110101011000111111111010010",
     496 => "00000110010010000111111111011000",  497 => "00000101111000110111111111011100",  498 => "00000101011111110111111111100001",  499 => "00000101000110110111111111100101",  500 => "00000100101101100111111111101001",  501 => "00000100010100100111111111101100",  502 => "00000011111011010111111111110000",  503 => "00000011100010010111111111110011",
     504 => "00000011001001000111111111110101",  505 => "00000010110000000111111111110111",  506 => "00000010010110110111111111111001",  507 => "00000001111101110111111111111011",  508 => "00000001100100100111111111111101",  509 => "00000001001011100111111111111110",  510 => "00000000110010010111111111111110",  511 => "00000000011001010111111111111111",
     512 => "00000000000000000111111111111111",  513 => "11111111100110110111111111111111",  514 => "11111111001101110111111111111110",  515 => "11111110110100100111111111111110",  516 => "11111110011011100111111111111101",  517 => "11111110000010010111111111111011",  518 => "11111101101001010111111111111001",  519 => "11111101010000000111111111110111",
     520 => "11111100110111000111111111110101",  521 => "11111100011101110111111111110011",  522 => "11111100000100110111111111110000",  523 => "11111011101011100111111111101100",  524 => "11111011010010100111111111101001",  525 => "11111010111001010111111111100101",  526 => "11111010100000010111111111100001",  527 => "11111010000111010111111111011100",
     528 => "11111001101110000111111111011000",  529 => "11111001010101000111111111010010",  530 => "11111000111011110111111111001101",  531 => "11111000100010110111111111000111",  532 => "11111000001001110111111111000001",  533 => "11110111110000100111111110111011",  534 => "11110111010111100111111110110100",  535 => "11110110111110100111111110101101",
     536 => "11110110100101100111111110100110",  537 => "11110110001100010111111110011111",  538 => "11110101110011010111111110010111",  539 => "11110101011010010111111110001111",  540 => "11110101000001010111111110000110",  541 => "11110100101000010111111101111101",  542 => "11110100001111000111111101110100",  543 => "11110011110110000111111101101011",
     544 => "11110011011101000111111101100001",  545 => "11110011000100000111111101010111",  546 => "11110010101011000111111101001101",  547 => "11110010010010000111111101000010",  548 => "11110001111001000111111100110111",  549 => "11110001100000000111111100101100",  550 => "11110001000111010111111100100001",  551 => "11110000101110010111111100010101",
     552 => "11110000010101010111111100001001",  553 => "11101111111100010111111011111100",  554 => "11101111100011100111111011101111",  555 => "11101111001010100111111011100010",  556 => "11101110110001100111111011010101",  557 => "11101110011000110111111011000111",  558 => "11101101111111110111111010111001",  559 => "11101101100111000111111010101011",
     560 => "11101101001110000111111010011100",  561 => "11101100110101010111111010001101",  562 => "11101100011100010111111001111110",  563 => "11101100000011100111111001101111",  564 => "11101011101010110111111001011111",  565 => "11101011010001110111111001001111",  566 => "11101010111001000111111000111110",  567 => "11101010100000010111111000101110",
     568 => "11101010000111100111111000011101",  569 => "11101001101110110111111000001011",  570 => "11101001010110000111110111111010",  571 => "11101000111101010111110111101000",  572 => "11101000100100100111110111010101",  573 => "11101000001100000111110111000011",  574 => "11100111110011010111110110110000",  575 => "11100111011010100111110110011101",
     576 => "11100111000001110111110110001001",  577 => "11100110101001010111110101110110",  578 => "11100110010000100111110101100010",  579 => "11100101111000000111110101001101",  580 => "11100101011111100111110100111001",  581 => "11100101000110110111110100100100",  582 => "11100100101110010111110100001110",  583 => "11100100010101110111110011111001",
     584 => "11100011111101010111110011100011",  585 => "11100011100100110111110011001101",  586 => "11100011001100010111110010110110",  587 => "11100010110011110111110010011111",  588 => "11100010011011010111110010001000",  589 => "11100010000010110111110001110001",  590 => "11100001101010010111110001011001",  591 => "11100001010010000111110001000001",
     592 => "11100000111001100111110000101001",  593 => "11100000100001010111110000010000",  594 => "11100000001000110111101111111000",  595 => "11011111110000100111101111011110",  596 => "11011111011000010111101111000101",  597 => "11011111000000000111101110101011",  598 => "11011110100111110111101110010001",  599 => "11011110001111100111101101110111",
     600 => "11011101110111010111101101011100",  601 => "11011101011111000111101101000001",  602 => "11011101000110110111101100100110",  603 => "11011100101110100111101100001010",  604 => "11011100010110100111101011101110",  605 => "11011011111110010111101011010010",  606 => "11011011100110010111101010110110",  607 => "11011011001110000111101010011001",
     608 => "11011010110110000111101001111100",  609 => "11011010011110000111101001011111",  610 => "11011010000110000111101001000001",  611 => "11011001101110000111101000100011",  612 => "11011001010110000111101000000101",  613 => "11011000111110000111100111100110",  614 => "11011000100110010111100111001000",  615 => "11011000001110010111100110101001",
     616 => "11010111110110100111100110001001",  617 => "11010111011110100111100101101010",  618 => "11010111000110110111100101001010",  619 => "11010110101111000111100100101001",  620 => "11010110010111010111100100001001",  621 => "11010101111111100111100011101000",  622 => "11010101100111110111100011000111",  623 => "11010101010000000111100010100101",
     624 => "11010100111000010111100010000100",  625 => "11010100100000110111100001100010",  626 => "11010100001001000111100000111111",  627 => "11010011110001100111100000011101",  628 => "11010011011001110111011111111010",  629 => "11010011000010010111011111010111",  630 => "11010010101010110111011110110011",  631 => "11010010010011010111011110001111",
     632 => "11010001111011110111011101101011",  633 => "11010001100100100111011101000111",  634 => "11010001001101000111011100100010",  635 => "11010000110101100111011011111110",  636 => "11010000011110010111011011011000",  637 => "11010000000111000111011010110011",  638 => "11001111101111110111011010001101",  639 => "11001111011000100111011001100111",
     640 => "11001111000001010111011001000001",  641 => "11001110101010000111011000011010",  642 => "11001110010010110111010111110011",  643 => "11001101111011110111010111001100",  644 => "11001101100100100111010110100101",  645 => "11001101001101100111010101111101",  646 => "11001100110110100111010101010101",  647 => "11001100011111010111010100101101",
     648 => "11001100001000010111010100000100",  649 => "11001011110001100111010011011011",  650 => "11001011011010100111010010110010",  651 => "11001011000011100111010010001000",  652 => "11001010101100110111010001011111",  653 => "11001010010110000111010000110101",  654 => "11001001111111000111010000001010",  655 => "11001001101000010111001111100000",
     656 => "11001001010001100111001110110101",  657 => "11001000111010110111001110001010",  658 => "11001000100100010111001101011110",  659 => "11001000001101100111001100110011",  660 => "11000111110111000111001100000111",  661 => "11000111100000100111001011011011",  662 => "11000111001001110111001010101110",  663 => "11000110110011010111001010000001",
     664 => "11000110011101000111001001010100",  665 => "11000110000110100111001000100111",  666 => "11000101110000000111000111111001",  667 => "11000101011001110111000111001011",  668 => "11000101000011100111000110011101",  669 => "11000100101101000111000101101111",  670 => "11000100010110110111000101000000",  671 => "11000100000000100111000100010001",
     672 => "11000011101010100111000011100010",  673 => "11000011010100010111000010110010",  674 => "11000010111110010111000010000011",  675 => "11000010101000000111000001010011",  676 => "11000010010010000111000000100010",  677 => "11000001111100000110111111110010",  678 => "11000001100110000110111111000001",  679 => "11000001010000010110111110010000",
     680 => "11000000111010010110111101011110",  681 => "11000000100100100110111100101100",  682 => "11000000001110110110111011111011",  683 => "10111111111000110110111011001000",  684 => "10111111100011010110111010010110",  685 => "10111111001101100110111001100011",  686 => "10111110110111110110111000110000",  687 => "10111110100010010110110111111101",
     688 => "10111110001100100110110111001001",  689 => "10111101110111000110110110010101",  690 => "10111101100001100110110101100001",  691 => "10111101001100000110110100101101",  692 => "10111100110110110110110011111000",  693 => "10111100100001010110110011000011",  694 => "10111100001100000110110010001110",  695 => "10111011110110110110110001011001",
     696 => "10111011100001100110110000100011",  697 => "10111011001100010110101111101101",  698 => "10111010110111000110101110110111",  699 => "10111010100010000110101110000001",  700 => "10111010001100110110101101001010",  701 => "10111001110111110110101100010011",  702 => "10111001100010110110101011011100",  703 => "10111001001101110110101010100100",
     704 => "10111000111001000110101001101101",  705 => "10111000100100000110101000110101",  706 => "10111000001111010110100111111101",  707 => "10110111111010100110100111000100",  708 => "10110111100101110110100110001011",  709 => "10110111010001000110100101010010",  710 => "10110110111100010110100100011001",  711 => "10110110100111110110100011100000",
     712 => "10110110010011000110100010100110",  713 => "10110101111110100110100001101100",  714 => "10110101101010000110100000110010",  715 => "10110101010101110110011111110111",  716 => "10110101000001010110011110111100",  717 => "10110100101101000110011110000001",  718 => "10110100011000110110011101000110",  719 => "10110100000100100110011100001010",
     720 => "10110011110000010110011011001111",  721 => "10110011011100000110011010010011",  722 => "10110011001000000110011001010110",  723 => "10110010110011110110011000011010",  724 => "10110010011111110110010111011101",  725 => "10110010001011110110010110100000",  726 => "10110001111000000110010101100011",  727 => "10110001100100000110010100100101",
     728 => "10110001010000010110010011101000",  729 => "10110000111100100110010010101010",  730 => "10110000101000110110010001101100",  731 => "10110000010101000110010000101101",  732 => "10110000000001010110001111101110",  733 => "10101111101101110110001110101111",  734 => "10101111011010010110001101110000",  735 => "10101111000110110110001100110001",
     736 => "10101110110011010110001011110001",  737 => "10101110011111110110001010110001",  738 => "10101110001100100110001001110001",  739 => "10101101111001010110001000110001",  740 => "10101101100110000110000111110000",  741 => "10101101010010110110000110101111",  742 => "10101100111111100110000101101110",  743 => "10101100101100100110000100101101",
     744 => "10101100011001010110000011101011",  745 => "10101100000110010110000010101010",  746 => "10101011110011100110000001101000",  747 => "10101011100000100110000000100101",  748 => "10101011001101110101111111100011",  749 => "10101010111010110101111110100000",  750 => "10101010101000000101111101011101",  751 => "10101010010101100101111100011010",
     752 => "10101010000010110101111011010111",  753 => "10101001110000010101111010010011",  754 => "10101001011101100101111001001111",  755 => "10101001001011010101111000001011",  756 => "10101000111000110101110111000111",  757 => "10101000100110010101110110000010",  758 => "10101000010100000101110100111110",  759 => "10101000000001110101110011111001",
     760 => "10100111101111100101110010110011",  761 => "10100111011101010101110001101110",  762 => "10100111001011010101110000101000",  763 => "10100110111001000101101111100010",  764 => "10100110100111000101101110011100",  765 => "10100110010101000101101101010110",  766 => "10100110000011010101101100001111",  767 => "10100101110001010101101011001001",
     768 => "10100101011111100101101010000010",  769 => "10100101001101110101101000111011",  770 => "10100100111100010101100111110011",  771 => "10100100101010100101100110101100",  772 => "10100100011001000101100101100100",  773 => "10100100000111100101100100011100",  774 => "10100011110110000101100011010011",  775 => "10100011100100100101100010001011",
     776 => "10100011010011010101100001000010",  777 => "10100011000001110101011111111001",  778 => "10100010110000100101011110110000",  779 => "10100010011111100101011101100111",  780 => "10100010001110010101011100011101",  781 => "10100001111101010101011011010011",  782 => "10100001101100010101011010001010",  783 => "10100001011011010101011000111111",
     784 => "10100001001010010101010111110101",  785 => "10100000111001100101010110101010",  786 => "10100000101000110101010101100000",  787 => "10100000011000000101010100010101",  788 => "10100000000111010101010011001001",  789 => "10011111110110110101010001111110",  790 => "10011111100110000101010000110010",  791 => "10011111010101100101001111100111",
     792 => "10011111000101010101001110011011",  793 => "10011110110100110101001101001110",  794 => "10011110100100100101001100000010",  795 => "10011110010100010101001010110101",  796 => "10011110000100000101001001101000",  797 => "10011101110011110101001000011011",  798 => "10011101100011110101000111001110",  799 => "10011101010011110101000110000001",
     800 => "10011101000011110101000100110011",  801 => "10011100110011110101000011100101",  802 => "10011100100100000101000010010111",  803 => "10011100010100010101000001001001",  804 => "10011100000100100100111111111011",  805 => "10011011110100110100111110101100",  806 => "10011011100101000100111101011101",  807 => "10011011010101100100111100001110",
     808 => "10011011000110000100111010111111",  809 => "10011010110110110100111001110000",  810 => "10011010100111010100111000100000",  811 => "10011010011000000100110111010001",  812 => "10011010001000110100110110000001",  813 => "10011001111001100100110100110001",  814 => "10011001101010100100110011100000",  815 => "10011001011011010100110010010000",
     816 => "10011001001100010100110000111111",  817 => "10011000111101100100101111101110",  818 => "10011000101110100100101110011101",  819 => "10011000011111110100101101001100",  820 => "10011000010001000100101011111011",  821 => "10011000000010010100101010101001",  822 => "10010111110011100100101001011000",  823 => "10010111100101000100101000000110",
     824 => "10010111010110100100100110110100",  825 => "10010111001000000100100101100001",  826 => "10010110111001110100100100001111",  827 => "10010110101011100100100010111100",  828 => "10010110011101010100100001101001",  829 => "10010110001111000100100000010110",  830 => "10010110000000110100011111000011",  831 => "10010101110010110100011101110000",
     832 => "10010101100100110100011100011100",  833 => "10010101010111000100011011001001",  834 => "10010101001001000100011001110101",  835 => "10010100111011010100011000100001",  836 => "10010100101101100100010111001101",  837 => "10010100011111110100010101111000",  838 => "10010100010010010100010100100100",  839 => "10010100000100110100010011001111",
     840 => "10010011110111010100010001111010",  841 => "10010011101001110100010000100101",  842 => "10010011011100100100001111010000",  843 => "10010011001111010100001101111011",  844 => "10010011000010000100001100100101",  845 => "10010010110100110100001011010000",  846 => "10010010100111110100001001111010",  847 => "10010010011010110100001000100100",
     848 => "10010010001101110100000111001110",  849 => "10010010000000110100000101110111",  850 => "10010001110100000100000100100001",  851 => "10010001100111010100000011001010",  852 => "10010001011010100100000001110011",  853 => "10010001001110000100000000011101",  854 => "10010001000001010011111111000101",  855 => "10010000110101000011111101101110",
     856 => "10010000101000100011111100010111",  857 => "10010000011100000011111010111111",  858 => "10010000001111110011111001101000",  859 => "10010000000011100011111000010000",  860 => "10001111110111100011110110111000",  861 => "10001111101011010011110101100000",  862 => "10001111011111010011110100000111",  863 => "10001111010011100011110010101111",
     864 => "10001111000111100011110001010110",  865 => "10001110111011110011101111111110",  866 => "10001110110000000011101110100101",  867 => "10001110100100010011101101001100",  868 => "10001110011000110011101011110010",  869 => "10001110001101010011101010011001",  870 => "10001110000001110011101001000000",  871 => "10001101110110010011100111100110",
     872 => "10001101101011000011100110001100",  873 => "10001101011111110011100100110011",  874 => "10001101010100100011100011011001",  875 => "10001101001001010011100001111110",  876 => "10001100111110010011100000100100",  877 => "10001100110011010011011111001010",  878 => "10001100101000100011011101101111",  879 => "10001100011101100011011100010101",
     880 => "10001100010010110011011010111010",  881 => "10001100001000000011011001011111",  882 => "10001011111101100011011000000100",  883 => "10001011110010110011010110101000",  884 => "10001011101000010011010101001101",  885 => "10001011011110000011010011110010",  886 => "10001011010011100011010010010110",  887 => "10001011001001010011010000111010",
     888 => "10001010111111000011001111011111",  889 => "10001010110100110011001110000011",  890 => "10001010101010110011001100100110",  891 => "10001010100000110011001011001010",  892 => "10001010010110110011001001101110",  893 => "10001010001101000011001000010001",  894 => "10001010000011010011000110110101",  895 => "10001001111001100011000101011000",
     896 => "10001001101111110011000011111011",  897 => "10001001100110010011000010011110",  898 => "10001001011100110011000001000001",  899 => "10001001010011010010111111100100",  900 => "10001001001010000010111110000111",  901 => "10001001000000100010111100101010",  902 => "10001000110111100010111011001100",  903 => "10001000101110010010111001101110",
     904 => "10001000100101010010111000010001",  905 => "10001000011100010010110110110011",  906 => "10001000010011010010110101010101",  907 => "10001000001010010010110011110111",  908 => "10001000000001100010110010011001",  909 => "10000111111000110010110000111010",  910 => "10000111110000010010101111011100",  911 => "10000111100111100010101101111101",
     912 => "10000111011111000010101100011111",  913 => "10000111010110110010101011000000",  914 => "10000111001110010010101001100001",  915 => "10000111000110000010101000000010",  916 => "10000110111101110010100110100011",  917 => "10000110110101110010100101000100",  918 => "10000110101101100010100011100101",  919 => "10000110100101100010100010000110",
     920 => "10000110011101110010100000100110",  921 => "10000110010101110010011111000111",  922 => "10000110001110000010011101100111",  923 => "10000110000110100010011100001000",  924 => "10000101111110110010011010101000",  925 => "10000101110111010010011001001000",  926 => "10000101101111110010010111101000",  927 => "10000101101000010010010110001000",
     928 => "10000101100001000010010100101000",  929 => "10000101011001110010010011001000",  930 => "10000101010010100010010001100111",  931 => "10000101001011100010010000000111",  932 => "10000101000100100010001110100110",  933 => "10000100111101100010001101000110",  934 => "10000100110110100010001011100101",  935 => "10000100101111110010001010000100",
     936 => "10000100101001000010001000100011",  937 => "10000100100010010010000111000010",  938 => "10000100011011110010000101100001",  939 => "10000100010101010010000100000000",  940 => "10000100001110110010000010011111",  941 => "10000100001000100010000000111110",  942 => "10000100000010000001111111011101",  943 => "10000011111100000001111101111011",
     944 => "10000011110101110001111100011010",  945 => "10000011101111110001111010111000",  946 => "10000011101001110001111001010111",  947 => "10000011100011110001110111110101",  948 => "10000011011110000001110110010011",  949 => "10000011011000010001110100110001",  950 => "10000011010010100001110011001111",  951 => "10000011001100110001110001101101",
     952 => "10000011000111010001110000001011",  953 => "10000011000001110001101110101001",  954 => "10000010111100100001101101000111",  955 => "10000010110111000001101011100101",  956 => "10000010110001110001101010000010",  957 => "10000010101100110001101000100000",  958 => "10000010100111100001100110111110",  959 => "10000010100010100001100101011011",
     960 => "10000010011101110001100011111001",  961 => "10000010011000110001100010010110",  962 => "10000010010100000001100000110011",  963 => "10000010001111010001011111010000",  964 => "10000010001010110001011101101110",  965 => "10000010000110000001011100001011",  966 => "10000010000001100001011010101000",  967 => "10000001111101010001011001000101",
     968 => "10000001111000110001010111100010",  969 => "10000001110100100001010101111111",  970 => "10000001110000100001010100011100",  971 => "10000001101100010001010010111001",  972 => "10000001101000010001010001010101",  973 => "10000001100100010001001111110010",  974 => "10000001100000100001001110001111",  975 => "10000001011100110001001100101011",
     976 => "10000001011001000001001011001000",  977 => "10000001010101010001001001100100",  978 => "10000001010001110001001000000001",  979 => "10000001001110010001000110011101",  980 => "10000001001010110001000100111010",  981 => "10000001000111100001000011010110",  982 => "10000001000100010001000001110010",  983 => "10000001000001000001000000001111",
     984 => "10000000111101110000111110101011",  985 => "10000000111010110000111101000111",  986 => "10000000110111110000111011100011",  987 => "10000000110101000000111010000000",  988 => "10000000110010010000111000011100",  989 => "10000000101111100000110110111000",  990 => "10000000101100110000110101010100",  991 => "10000000101010010000110011110000",
     992 => "10000000100111110000110010001100",  993 => "10000000100101010000110000101000",  994 => "10000000100011000000101111000100",  995 => "10000000100000110000101101011111",  996 => "10000000011110100000101011111011",  997 => "10000000011100010000101010010111",  998 => "10000000011010010000101000110011",  999 => "10000000011000010000100111001111",
    1000 => "10000000010110100000100101101010", 1001 => "10000000010100110000100100000110", 1002 => "10000000010011000000100010100010", 1003 => "10000000010001010000100000111110", 1004 => "10000000001111110000011111011001", 1005 => "10000000001110010000011101110101", 1006 => "10000000001100110000011100010001", 1007 => "10000000001011100000011010101100",
    1008 => "10000000001010000000011001001000", 1009 => "10000000001001000000010111100011", 1010 => "10000000000111110000010101111111", 1011 => "10000000000110110000010100011011", 1012 => "10000000000101110000010010110110", 1013 => "10000000000101000000010001010010", 1014 => "10000000000100000000001111101101", 1015 => "10000000000011010000001110001001",
    1016 => "10000000000010110000001100100100", 1017 => "10000000000010010000001011000000", 1018 => "10000000000001110000001001011011", 1019 => "10000000000001010000000111110111", 1020 => "10000000000000110000000110010010", 1021 => "10000000000000100000000100101110", 1022 => "10000000000000100000000011001001", 1023 => "10000000000000010000000001100101"
  );

  signal m_lut          : std_logic_vector_array_t(2 ** DDS_SIN_LOOKUP_INDEX_WIDTH - 1 downto 0)(LUT_WIDTH - 1 downto 0) := LUT_INIT;

  signal r0_read_half   : std_logic;
  signal r0_read_data   : std_logic_vector(LUT_WIDTH - 1 downto 0);

  signal r1_read_half   : std_logic;
  signal r1_read_data   : std_logic_vector(LUT_WIDTH - 1 downto 0);
  signal w1_data_i      : signed(LUT_WIDTH/2 - 1 downto 0);
  signal w1_data_q      : signed(LUT_WIDTH/2 - 1 downto 0);
  signal w1_data_i_inv  : signed(LUT_WIDTH/2 - 1 downto 0);
  signal w1_data_q_inv  : signed(LUT_WIDTH/2 - 1 downto 0);

begin

  assert (LATENCY = 3)
    report "LATENCY expected to be 3"
    severity failure;

  assert (DATA_WIDTH = LUT_WIDTH/2)
    report "DATA_WIDTH must be = LUT_WIDTH/2, otherwise max negative->invert behavior is not guaranteed"
    severity failure;

  process(Clk)
  begin
    if rising_edge(Clk) then
      r0_read_half <= Read_half;
      r0_read_data <= m_lut(to_integer(Read_index));
    end if;
  end process;

  process(Clk)
  begin
    if rising_edge(Clk) then
      r1_read_half <= r0_read_half;
      r1_read_data <= r0_read_data;
    end if;
  end process;

  (w1_data_q, w1_data_i) <= signed(r1_read_data);
  w1_data_i_inv <= -w1_data_i;
  w1_data_q_inv <= -w1_data_q;

  -- PSL underflow_i : assert always (w1_data_i(LUT_WIDTH/2 - 1) = '1') -> (or_reduce(w1_data_i(LUT_WIDTH/2 - 2 downto 0)) = '1');
  -- PSL underflow_q : assert always (w1_data_q(LUT_WIDTH/2 - 1) = '1') -> (or_reduce(w1_data_q(LUT_WIDTH/2 - 2 downto 0)) = '1');

  process(Clk)
  begin
    if rising_edge(Clk) then
      if (r1_read_half = '0') then
        Read_data(0) <= w1_data_i(LUT_WIDTH/2 - 1 downto (LUT_WIDTH/2 - DATA_WIDTH));
        Read_data(1) <= w1_data_q(LUT_WIDTH/2 - 1 downto (LUT_WIDTH/2 - DATA_WIDTH));
      else
        Read_data(0) <= w1_data_i_inv(LUT_WIDTH/2 - 1 downto (LUT_WIDTH/2 - DATA_WIDTH));
        Read_data(1) <= w1_data_q_inv(LUT_WIDTH/2 - 1 downto (LUT_WIDTH/2 - DATA_WIDTH));
      end if;
    end if;
  end process;

end architecture rtl;
