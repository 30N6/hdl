library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library common_lib;
  use common_lib.common_pkg.all;
  use common_lib.math_pkg.all;

library dsp_lib;
  use dsp_lib.dsp_pkg.all;

entity synthesizer_16 is
generic (
  INPUT_DATA_WIDTH  : natural;
  OUTPUT_DATA_WIDTH : natural
);
port (
  Clk                       : in  std_logic;
  Rst                       : in  std_logic;

  Input_ctrl                : in  synthesizer_control_t;
  Input_data                : in  signed_array_t(1 downto 0)(INPUT_DATA_WIDTH - 1 downto 0);

  Output_valid              : out std_logic;
  Output_data               : out signed_array_t(1 downto 0)(OUTPUT_DATA_WIDTH - 1 downto 0);

  Error_stretcher_overflow  : out std_logic;
  Error_stretcher_underflow : out std_logic;
  Error_filter_overflow     : out std_logic;
  Error_mux_input_overflow  : out std_logic;
  Error_mux_fifo_overflow   : out std_logic;
  Error_mux_fifo_underflow  : out std_logic
);
end entity synthesizer_16;

architecture rtl of synthesizer_16 is

  constant NUM_CHANNELS : natural := 16;
  constant NUM_COEFS    : natural := 128;
  constant COEF_WIDTH   : natural := 20;
  constant COEF_DATA    : signed_array_t(NUM_COEFS - 1 downto 0)(COEF_WIDTH - 1 downto 0) := (
      0 => "00000000000001101011",   1 => "00000000000000100000",   2 => "11111111111110010011",   3 => "11111111111010111000",   4 => "11111111110110001011",   5 => "11111111110000001100",   6 => "11111111101001000101",   7 => "11111111100001001000",
      8 => "11111111011000110101",   9 => "11111111010000110001",  10 => "11111111001001101110",  11 => "11111111000100100110",  12 => "11111111000010010110",  13 => "11111111000011111100",  14 => "11111111001010010101",  15 => "11111111010110010100",
     16 => "11111111101000011110",  17 => "00000000000001000111",  18 => "00000000100000001000",  19 => "00000001000100111111",  20 => "00000001101110101000",  21 => "00000010011011100000",  22 => "00000011001001100001",  23 => "00000011110110000111",
     24 => "00000100011110010011",  25 => "00000100111110110101",  26 => "00000101010100010000",  27 => "00000101011011001110",  28 => "00000101010000100101",  29 => "00000100110001101001",  30 => "00000011111100011010",  31 => "00000010101111110010",
     32 => "00000001001011110000",  33 => "11111111010001101000",  34 => "11111101000100000100",  35 => "11111010100111001011",  36 => "11111000000000100100",  37 => "11110101010111001100",  38 => "11110010110011001111",  39 => "11110000011101111001",
     40 => "11101110100001000011",  41 => "11101101000110111011",  42 => "11101100011001101011",  43 => "11101100100010111011",  44 => "11101101101011010101",  45 => "11101111111010000111",  46 => "11110011010100101001",  47 => "11110111111110000011",
     48 => "11111101110110111010",  49 => "00000100111101000011",  50 => "00001101001011011101",  51 => "00010110011010001111",  52 => "00100000011110110000",  53 => "00101011001011111000",  54 => "00110110010010010111",  55 => "01000001100001010000",
     56 => "01001100100110011111",  57 => "01010111001111100000",  58 => "01100001001001110110",  59 => "01101010000011111010",  60 => "01110001101101100000",  61 => "01110111111000100010",  62 => "01111100011001011101",  63 => "01111111000111110100",
     64 => "01111111111110100001",  65 => "01111110111011111110",  66 => "01111100000010010010",  67 => "01110111010111000001",  68 => "01110001000011001000",  69 => "01101001010010011111",  70 => "01100000010011100000",  71 => "01010110010110100001",
     72 => "01001011101101010000",  73 => "01000000101010000111",  74 => "00110101011111100001",  75 => "00101010011111010100",  76 => "00011111111010001000",  77 => "00010101111110110011",  78 => "00001100111010000010",  79 => "00000100110110000001",
     80 => "11111101111010001010",  81 => "11111000001011000011",  82 => "11110011101010011101",  83 => "11110000010111011100",  84 => "11101110001110100111",  85 => "11101101001010011011",  86 => "11101101000011100100",  87 => "11101101110001010110",
     88 => "11101111001010001110",  89 => "11110001000100001110",  90 => "11110011010101010011",  91 => "11110101110011111000",  92 => "11111000010111000100",  93 => "11111010110110111111",  94 => "11111101001101000010",  95 => "11111111010011111100",
     96 => "00000001000111110101",  97 => "00000010100110010100",  98 => "00000011101110010001",  99 => "00000100011111110111", 100 => "00000100111100001111", 101 => "00000101000101011010", 102 => "00000100111110000100", 103 => "00000100101001001110",
    104 => "00000100001010001010", 105 => "00000011100100001000", 106 => "00000010111010001110", 107 => "00000010001111001111", 108 => "00000001100101100011", 109 => "00000000111111000110", 110 => "00000000011101010010", 111 => "00000000000001000000",
    112 => "11111111101010101111", 113 => "11111111011010100000", 114 => "11111111001111111101", 115 => "11111111001010100010", 116 => "11111111001001011100", 117 => "11111111001011110001", 118 => "11111111010000101000", 119 => "11111111010111000110",
    120 => "11111111011110011000", 121 => "11111111100101110010", 122 => "11111111101100110001", 123 => "11111111110010111011", 124 => "11111111111000000001", 125 => "11111111111011111011", 126 => "11111111111110101100", 127 => "00000000000000011000"
  );

begin

  i_synthesizer : entity dsp_lib.synthesizer_common
  generic map (
    INPUT_DATA_WIDTH  => INPUT_DATA_WIDTH,
    OUTPUT_DATA_WIDTH => OUTPUT_DATA_WIDTH,
    NUM_CHANNELS      => NUM_CHANNELS,
    NUM_COEFS         => NUM_COEFS,
    COEF_WIDTH        => COEF_WIDTH,
    COEF_DATA         => COEF_DATA
  )
  port map (
    Clk                       => Clk,
    Rst                       => Rst,


    Input_ctrl                => Input_ctrl,
    Input_data                => Input_data,

    Output_valid              => Output_valid,
    Output_data               => Output_data,

    Error_stretcher_overflow  => Error_stretcher_overflow,
    Error_stretcher_underflow => Error_stretcher_underflow,
    Error_filter_overflow     => Error_filter_overflow,
    Error_mux_input_overflow  => Error_mux_input_overflow,
    Error_mux_fifo_overflow   => Error_mux_fifo_overflow,
    Error_mux_fifo_underflow  => Error_mux_fifo_underflow
  );

end architecture rtl;
